module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49,  o);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49;
output o;
wire x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31_c, x32_c, x33_c, x34_c, x35_c, x36_c, x37_c, x38_c, x39_c, x40_c, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49_c;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49;
assign x0_c = ~x0;
assign x1_c = ~x1;
assign x2_c = ~x2;
assign x3_c = ~x3;
assign x4_c = ~x4;
assign x5_c = ~x5;
assign x6_c = ~x6;
assign x7_c = ~x7;
assign x8_c = ~x8;
assign x9_c = ~x9;
assign x10_c = ~x10;
assign x11_c = ~x11;
assign x12_c = ~x12;
assign x13_c = ~x13;
assign x14_c = ~x14;
assign x15_c = ~x15;
assign x16_c = ~x16;
assign x17_c = ~x17;
assign x18_c = ~x18;
assign x19_c = ~x19;
assign x20_c = ~x20;
assign x21_c = ~x21;
assign x22_c = ~x22;
assign x23_c = ~x23;
assign x24_c = ~x24;
assign x25_c = ~x25;
assign x26_c = ~x26;
assign x27_c = ~x27;
assign x28_c = ~x28;
assign x29_c = ~x29;
assign x30_c = ~x30;
assign x31_c = ~x31;
assign x32_c = ~x32;
assign x33_c = ~x33;
assign x34_c = ~x34;
assign x35_c = ~x35;
assign x36_c = ~x36;
assign x37_c = ~x37;
assign x38_c = ~x38;
assign x39_c = ~x39;
assign x40_c = ~x40;
assign x41_c = ~x41;
assign x42_c = ~x42;
assign x43_c = ~x43;
assign x44_c = ~x44;
assign x45_c = ~x45;
assign x46_c = ~x46;
assign x47_c = ~x47;
assign x48_c = ~x48;
assign x49_c = ~x49;
and (w0, x0, x1, x4_c, x5, x6, x8_c, x10, x11_c, x12, x13_c, x15_c, x16_c, x17_c, x20_c, x21_c, x22, x26, x28_c, x29_c, x32_c, x33, x34, x35_c, x36, x38, x39_c, x41, x42, x45, x47_c, x48);
and (w1, x2_c, x4_c, x20_c, x25, x29_c);
and (w2, x11_c, x15_c, x17_c, x22, x24, x25_c, x33_c, x35, x39_c, x42_c, x45_c);
and (w3, x1_c, x2_c, x4_c, x9, x10_c, x11, x15, x16, x17_c, x20_c, x21_c, x22, x24, x26_c, x28_c, x30, x32, x34_c, x35, x36, x38, x39_c, x43_c, x44, x46, x47_c, x49_c);
and (w4, x6, x8, x10, x12_c, x15_c, x18, x24_c, x25, x28, x29, x31, x34_c, x38, x39_c, x42, x45, x46_c, x48_c, x49);
and (w5, x0, x2_c, x3_c, x4, x13_c, x15, x17_c, x19, x20_c, x24, x25, x28_c, x29, x33, x35_c, x40_c, x43_c, x44_c, x46, x47);
and (w6, x4, x7_c, x9_c, x10_c, x16, x17_c, x26_c, x33_c, x35_c, x38, x40, x48_c);
and (w7, x2, x3, x4_c, x5, x7_c, x8, x9_c, x12, x13, x17, x19, x20, x23, x24, x30, x32_c, x34, x35, x38_c, x40, x41, x42, x43_c, x46);
and (w8, x0, x2_c, x3_c, x4, x5, x6, x8_c, x9_c, x12, x17, x18_c, x19_c, x24, x25_c, x26_c, x28, x29_c, x31, x32_c, x33, x36, x37_c, x38, x39_c, x41_c, x44, x45, x48_c, x49);
and (w9, x3_c, x15_c, x16_c, x17, x18_c, x31, x32_c, x36, x41, x48);
and (w10, x39, x43_c, x45);
and (w11, x0, x1, x2_c, x3, x4_c, x5, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14_c, x15_c, x16, x17, x18, x19, x20, x21, x22, x23_c, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33, x34_c, x35_c, x36_c, x37, x38, x39, x40_c, x42_c, x43_c, x44_c, x45_c, x46, x47, x48, x49);
and (w12, x0, x1, x2_c, x3, x4_c, x5_c, x7_c, x8_c, x9_c, x10, x11, x12_c, x13_c, x14, x16, x17_c, x18_c, x19_c, x20, x21, x22_c, x23_c, x27_c, x29_c, x31_c, x32_c, x33_c, x35_c, x36, x37, x39, x40, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48, x49_c);
and (w13, x15_c, x21, x44_c, x47);
and (w14, x0, x2_c, x3, x5, x7, x10, x12, x13, x15, x17, x21_c, x24_c, x26_c, x27_c, x31, x32, x34_c, x39_c, x41, x42, x45_c, x46_c, x49);
and (w15, x0_c, x1, x2, x3, x4, x5_c, x6_c, x7_c, x8_c, x10, x12_c, x13_c, x14, x15, x16_c, x18, x19_c, x20_c, x21_c, x22_c, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x32_c, x33, x34_c, x35, x36, x37_c, x38, x40, x41, x43, x44, x45_c, x46, x47, x48_c, x49);
and (w16, x14, x15, x26, x27_c, x31_c, x35, x38, x42_c, x45_c, x46_c, x48);
and (w17, x1, x3, x11, x14_c, x20_c, x21_c, x31_c, x40_c, x43_c, x45_c, x46, x47_c);
and (w18, x1, x6, x8_c, x9, x22, x26_c, x27, x28_c, x30_c, x36, x38, x39_c, x42, x44_c, x47_c, x49);
and (w19, x0, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9, x13, x14_c, x15, x16, x17, x18_c, x19, x20_c, x21_c, x22_c, x24, x25, x26_c, x27_c, x28_c, x29, x30_c, x31_c, x33_c, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41_c, x42_c, x43_c, x44_c, x45, x47, x48, x49_c);
and (w20, x0_c, x1_c, x4_c, x5_c, x6_c, x7_c, x9_c, x10, x15_c, x16, x22_c, x24_c, x25_c, x27_c, x28, x30_c, x31_c, x32, x34, x35, x37, x38, x41_c, x42_c, x44, x48, x49);
and (w21, x4, x5_c, x7_c, x9_c, x10_c, x12, x16, x18, x19_c, x20_c, x22, x24_c, x26, x27, x30, x38_c, x43_c, x45, x48);
and (w22, x0, x3, x4, x6, x11_c, x14, x16, x17, x20, x21, x23_c, x26, x27_c, x28_c, x29_c, x30_c, x34_c, x36, x43_c);
and (w23, x0, x4_c, x7, x8_c, x9_c, x13_c, x16, x18_c, x21, x23, x25_c, x27_c, x28_c, x29_c, x32, x34_c, x37, x39, x40_c, x41, x45, x47, x48_c, x49_c);
and (w24, x0_c, x2_c, x4, x9_c, x11, x12, x14_c, x15, x18_c, x24, x28, x29, x32, x33, x34, x37, x38_c, x40_c, x47);
and (w25, x0, x1_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23, x24, x25_c, x26_c, x27_c, x29, x30, x32, x33_c, x35_c, x36, x37_c, x38_c, x39, x40_c, x41_c, x42, x43_c, x44, x45, x46, x47_c, x48);
and (w26, x0_c, x1, x2, x3_c, x4_c, x5, x6_c, x7_c, x8, x9_c, x10, x12_c, x14_c, x15_c, x16, x17, x20_c, x22_c, x24, x25_c, x27_c, x28, x29, x30_c, x31, x33, x34_c, x35, x36_c, x37_c, x38_c, x39, x40, x41_c, x42_c, x43, x44_c, x45, x46, x47, x49);
and (w27, x0, x1_c, x2, x4, x5, x6, x7_c, x8_c, x9, x10, x11, x12, x14, x17_c, x19_c, x20_c, x21_c, x22_c, x23, x25_c, x26_c, x27, x28, x29, x33_c, x34, x37_c, x39_c, x41_c, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c);
and (w28, x0_c, x1, x2, x3_c, x4_c, x5, x6, x7_c, x8_c, x9_c, x10, x11_c, x12, x13_c, x14_c, x17_c, x18_c, x19, x20, x23, x24_c, x26, x27_c, x28_c, x29_c, x30, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x38_c, x39, x40, x41, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c);
assign w29 = x48;
and (w30, x1_c, x4, x6, x9, x13, x14_c, x17, x21, x22_c, x26_c, x27, x28_c, x32, x34_c, x38, x41_c, x45_c, x46, x47, x48);
and (w31, x0_c, x1_c, x6_c, x7, x10_c, x11, x23_c, x25_c, x36_c, x40_c, x43, x47, x48_c);
and (w32, x0, x1_c, x2, x3_c, x4, x5, x6, x7, x8_c, x9_c, x10, x11, x12_c, x13, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20, x23, x24, x25_c, x26_c, x27_c, x28_c, x29, x30, x31_c, x32_c, x33, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x44, x45_c, x46_c, x47, x48_c);
and (w33, x0_c, x1, x3, x5, x11_c, x12, x13_c, x14_c, x15_c, x17, x18_c, x19_c, x20_c, x22, x23_c, x24, x25, x26_c, x27, x28, x29, x31, x32_c, x33, x34_c, x36_c, x37_c, x38_c, x39, x40, x42_c, x43, x44_c, x45, x46_c, x47, x48_c, x49);
and (w34, x0_c, x2, x4, x8_c, x10_c, x12_c, x13, x14_c, x17, x19_c, x21_c, x23_c, x24, x25_c, x26, x28_c, x30_c, x32_c, x34, x35, x37_c, x38_c, x39, x40_c, x41, x43_c, x44_c, x45, x47, x48, x49_c);
and (w35, x0, x1_c, x2, x3_c, x4_c, x5, x6, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14_c, x15, x16, x17, x18, x19_c, x20, x21, x22, x23, x24, x25, x26, x27_c, x28, x29, x30_c, x31_c, x32, x33_c, x34_c, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42, x43, x44_c, x45_c, x46_c, x47, x48_c, x49_c);
and (w36, x4, x5, x17, x18, x19_c, x22, x35_c, x38_c, x42, x43_c, x44_c);
assign w37 = x16_c;
and (w38, x0_c, x6, x7, x9, x12_c, x13, x14_c, x16_c, x17_c, x20, x21, x22, x23, x24, x25_c, x28, x29, x34_c, x36_c, x37, x38, x39_c, x40_c, x42_c, x43, x46_c, x48_c);
and (w39, x0, x1_c, x3_c, x4_c, x6_c, x7, x9_c, x13, x16_c, x20_c, x23_c, x25_c, x26_c, x27, x28_c, x30, x31_c, x32_c, x34_c, x35, x36, x37_c, x38, x40_c, x41, x42_c, x45_c, x46_c, x47, x48_c, x49);
and (w40, x1, x3, x4, x5, x6_c, x12, x14_c, x15_c, x18, x19_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x32, x34, x35_c, x38, x49);
and (w41, x0, x1_c, x2_c, x3_c, x6_c, x7_c, x9_c, x10, x12_c, x13, x14, x16, x17, x18_c, x22, x23_c, x32_c, x33_c, x34, x38, x39_c, x40, x41, x42, x43_c, x44_c, x46, x47, x48, x49_c);
and (w42, x3, x9, x16_c, x20, x23, x31_c, x32_c, x33_c, x36_c, x41, x44, x48_c);
and (w43, x0_c, x2_c, x3_c, x5, x6, x7, x8, x9, x11_c, x12, x13_c, x15_c, x18, x19, x21, x22_c, x23_c, x24_c, x25_c, x28_c, x29, x30, x32, x33_c, x34_c, x38, x39, x42, x43_c, x45, x46, x47_c, x48_c);
and (w44, x10, x19_c, x35_c);
and (w45, x1, x2_c, x3_c, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x11, x12, x13_c, x14_c, x15, x16, x17, x18, x19, x20_c, x21, x22_c, x23_c, x24_c, x25_c, x26_c, x27, x28, x29, x30_c, x31_c, x32_c, x33_c, x34, x35, x36_c, x37_c, x38, x39_c, x40, x41, x43_c, x44_c, x45, x46_c, x47, x48_c, x49_c);
and (w46, x0, x1, x2_c, x3_c, x5, x6, x7_c, x10, x11_c, x12, x13, x16_c, x23, x24, x33, x36, x37_c, x38, x43_c, x44, x46, x49);
and (w47, x2_c, x3, x6, x10, x12, x14, x21_c, x22, x26, x27_c, x31_c, x32, x34_c, x40, x41_c, x43_c, x44, x47_c, x49);
and (w48, x1_c, x18, x23, x31, x32_c, x33, x36, x48_c);
and (w49, x0_c, x1, x2_c, x3_c, x4_c, x6, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14_c, x15, x16_c, x17_c, x18, x19_c, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x27, x29_c, x30, x31_c, x32, x34, x35_c, x36, x38_c, x39_c, x40, x41_c, x42_c, x43, x44_c, x45, x46, x47, x48, x49);
xor (o, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49);
endmodule
