module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99,  o);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99;
output o;
wire x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31_c, x32_c, x33_c, x34_c, x35_c, x36_c, x37_c, x38_c, x39_c, x40_c, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98_c, x99_c;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757;
assign x0_c = ~x0;
assign x1_c = ~x1;
assign x2_c = ~x2;
assign x3_c = ~x3;
assign x4_c = ~x4;
assign x5_c = ~x5;
assign x6_c = ~x6;
assign x7_c = ~x7;
assign x8_c = ~x8;
assign x9_c = ~x9;
assign x10_c = ~x10;
assign x11_c = ~x11;
assign x12_c = ~x12;
assign x13_c = ~x13;
assign x14_c = ~x14;
assign x15_c = ~x15;
assign x16_c = ~x16;
assign x17_c = ~x17;
assign x18_c = ~x18;
assign x19_c = ~x19;
assign x20_c = ~x20;
assign x21_c = ~x21;
assign x22_c = ~x22;
assign x23_c = ~x23;
assign x24_c = ~x24;
assign x25_c = ~x25;
assign x26_c = ~x26;
assign x27_c = ~x27;
assign x28_c = ~x28;
assign x29_c = ~x29;
assign x30_c = ~x30;
assign x31_c = ~x31;
assign x32_c = ~x32;
assign x33_c = ~x33;
assign x34_c = ~x34;
assign x35_c = ~x35;
assign x36_c = ~x36;
assign x37_c = ~x37;
assign x38_c = ~x38;
assign x39_c = ~x39;
assign x40_c = ~x40;
assign x41_c = ~x41;
assign x42_c = ~x42;
assign x43_c = ~x43;
assign x44_c = ~x44;
assign x45_c = ~x45;
assign x46_c = ~x46;
assign x47_c = ~x47;
assign x48_c = ~x48;
assign x49_c = ~x49;
assign x50_c = ~x50;
assign x51_c = ~x51;
assign x52_c = ~x52;
assign x53_c = ~x53;
assign x54_c = ~x54;
assign x55_c = ~x55;
assign x56_c = ~x56;
assign x57_c = ~x57;
assign x58_c = ~x58;
assign x59_c = ~x59;
assign x60_c = ~x60;
assign x61_c = ~x61;
assign x62_c = ~x62;
assign x63_c = ~x63;
assign x64_c = ~x64;
assign x65_c = ~x65;
assign x66_c = ~x66;
assign x67_c = ~x67;
assign x68_c = ~x68;
assign x69_c = ~x69;
assign x70_c = ~x70;
assign x71_c = ~x71;
assign x72_c = ~x72;
assign x73_c = ~x73;
assign x74_c = ~x74;
assign x75_c = ~x75;
assign x76_c = ~x76;
assign x77_c = ~x77;
assign x78_c = ~x78;
assign x79_c = ~x79;
assign x80_c = ~x80;
assign x81_c = ~x81;
assign x82_c = ~x82;
assign x83_c = ~x83;
assign x84_c = ~x84;
assign x85_c = ~x85;
assign x86_c = ~x86;
assign x87_c = ~x87;
assign x88_c = ~x88;
assign x89_c = ~x89;
assign x90_c = ~x90;
assign x91_c = ~x91;
assign x92_c = ~x92;
assign x93_c = ~x93;
assign x94_c = ~x94;
assign x95_c = ~x95;
assign x96_c = ~x96;
assign x97_c = ~x97;
assign x98_c = ~x98;
assign x99_c = ~x99;
and (w0, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92_c, x93_c, x95_c, x96, x98, x99);
and (w1, x24, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2, x3_c, x10_c, x14_c, x21_c, x29, x34_c, x41_c, x43, x81, x84_c, x86, x99_c);
and (w3, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x37, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x77_c, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x77_c, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w7, x2_c, x3, x4_c, x5, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w8, x2_c, x6_c, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w9, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w10, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w11, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x38_c, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w12, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x47, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w13, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x20, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w14, x16, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w15, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92, x96, x97_c);
and (w16, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w17, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x44_c, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w18, x0_c, x4, x17, x57, x75_c, x83, x90_c);
and (w19, x0_c, x5, x23_c, x30_c, x31_c, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w20, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82_c, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w21, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w22, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w23, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w24, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w25, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x56_c, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w26, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w27, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w28, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35_c, x83_c);
and (w29, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x15_c, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w30, x13_c, x14_c, x37_c, x39_c, x45_c, x53, x82, x90_c, x96, x98, x99_c);
and (w31, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x56_c, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w32, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x66_c, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w33, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w34, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x90, x91_c, x95, x96, x97, x99_c);
and (w35, x1_c, x3_c, x9, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w36, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w37, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w38, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w39, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x53_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w40, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82, x83_c);
and (w41, x0_c, x1, x2_c, x3, x4, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25, x26, x27_c, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36_c, x37_c, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48, x49, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57_c, x58, x59, x60, x61, x62, x63_c, x64_c, x65_c, x66, x67, x68_c, x69, x70_c, x71, x72, x73, x74, x75_c, x76, x77, x78, x79_c, x80_c, x81, x82_c, x83, x84, x85, x86, x87_c, x88_c, x89, x90_c, x92_c, x93_c, x94, x95, x96, x97, x98, x99);
and (w42, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x46, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w43, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w44, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x47, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w45, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w46, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x77, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w47, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w48, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w49, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x50_c, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w50, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x14, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w51, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x23, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w52, x0, x2, x7_c, x8, x15_c, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w53, x12_c, x32, x86_c, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w54, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w55, x0_c, x2, x3, x4_c, x7, x8, x11, x15_c, x16_c, x17_c, x18, x22, x24, x26_c, x28_c, x30, x31_c, x32, x34_c, x35_c, x36, x37, x38_c, x40, x41, x42_c, x44, x45, x46, x47, x48, x49_c, x53_c, x54, x56_c, x57, x58_c, x60, x61, x62_c, x63, x64, x65_c, x66_c, x67_c, x68_c, x70_c, x72_c, x73, x75, x76_c, x77, x78, x81_c, x82, x83, x85_c, x88, x90, x91, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w56, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w57, x3, x5_c, x6, x7, x8_c, x13, x15_c, x16_c, x18_c, x19, x21, x22_c, x26, x28, x31, x33_c, x34, x38, x39_c, x42_c, x47_c, x48_c, x49_c, x50_c, x51, x53, x54, x56_c, x57, x58_c, x59_c, x62, x63, x66_c, x69_c, x70_c, x73, x74_c, x75, x76_c, x81, x83_c, x84, x87, x89_c, x90_c, x93_c, x94_c, x96, x99_c);
and (w58, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71, x72_c, x81, x84, x85, x95, x99);
and (w59, x0, x1_c, x2, x3_c, x4, x5_c, x6_c, x7_c, x9, x10, x11, x13_c, x15, x16, x17_c, x18, x19, x21, x22, x23, x24, x25_c, x26_c, x27, x30, x31_c, x33, x34_c, x36_c, x37, x38, x39_c, x40_c, x42, x43, x44, x45_c, x46, x47_c, x48, x49_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x59_c, x60_c, x61, x62, x63, x64, x65, x66, x68_c, x69, x71, x72_c, x73_c, x74_c, x76_c, x77_c, x79, x80, x81, x82, x86_c, x88_c, x89_c, x90, x91_c, x92, x93_c, x96_c, x98_c, x99_c);
and (w60, x11_c, x13, x15_c, x18_c, x22_c, x26_c, x27_c, x30_c, x36, x37_c, x39, x42_c, x45, x50, x51_c, x54_c, x56, x60, x63_c, x66_c, x71_c, x72, x81, x85_c, x90_c, x97_c, x98_c);
and (w61, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w62, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25_c, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w63, x26, x33_c, x44, x53);
and (w64, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w65, x2_c, x12, x16_c, x17_c, x18_c, x25, x29, x34_c, x40_c, x41_c, x44, x46_c, x50_c, x51_c, x53_c, x56, x58_c, x59, x60, x61_c, x65_c, x66_c, x71_c, x80_c, x82_c, x83, x84, x87, x91_c, x93_c, x95_c, x96_c);
and (w66, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w67, x1, x2_c, x7, x9_c, x10_c, x12, x13_c, x14, x15_c, x16_c, x18, x19, x21, x23_c, x27_c, x29_c, x31_c, x33_c, x34, x35, x38_c, x41_c, x42, x45, x46_c, x47_c, x48_c, x50, x52, x53_c, x56, x58_c, x59_c, x60, x62_c, x63, x64, x66_c, x69_c, x70_c, x71_c, x74, x75, x76, x78, x79_c, x86, x87_c, x88_c, x89, x90, x91_c, x92, x93, x94, x95, x96, x97);
and (w68, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w69, x1, x2_c, x3, x4, x5, x8_c, x9, x11_c, x12, x13, x15_c, x17, x18, x19, x21, x22_c, x23_c, x25, x29_c, x34, x37, x38_c, x39_c, x40, x41_c, x43_c, x45, x46_c, x49_c, x52, x53, x55_c, x56_c, x57, x58, x60, x61_c, x64_c, x69, x72, x74_c, x76, x77, x79, x80_c, x84, x86, x87, x88, x89, x91, x92, x93, x94, x96, x97, x98, x99_c);
and (w70, x2_c, x11, x26, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w71, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x32_c, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w72, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x56, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w73, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50, x82, x90_c, x96, x98, x99_c);
and (w74, x7, x13, x14, x15_c, x35_c, x37_c, x60, x70, x79, x88, x93_c);
and (w75, x12_c, x32, x71_c, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w76, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w77, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x50, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w78, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x81, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w79, x4_c, x10, x15_c, x22_c, x24_c, x27_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w80, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w81, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x66_c, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w82, x0, x3, x4, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w83, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x78, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w84, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88, x91_c, x92_c, x93_c, x96, x97_c);
and (w85, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x18_c, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w86, x1_c, x3_c, x4_c, x5_c, x6, x9_c, x10, x11_c, x13, x17, x20, x22_c, x23, x25_c, x26_c, x28, x29_c, x30_c, x31, x35, x37_c, x40, x42_c, x43_c, x49, x51, x52_c, x53, x54, x57_c, x58_c, x59_c, x61, x62_c, x64, x66, x67_c, x69, x70, x71, x72_c, x73, x75, x80_c, x81_c, x85, x86_c, x88_c, x89, x93_c, x95_c, x96, x98_c, x99_c);
and (w87, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x66_c, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w88, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w89, x0_c, x2_c, x3_c, x6, x7_c, x10, x11, x14_c, x15_c, x16, x17, x21_c, x23_c, x25, x27, x28_c, x29, x30, x31_c, x32, x35_c, x36, x38, x39, x41_c, x42, x43_c, x44_c, x45_c, x46, x49_c, x52_c, x54_c, x57, x58, x59, x61, x65, x66_c, x67_c, x70, x71_c, x72_c, x74_c, x75, x76_c, x78_c, x79_c, x80_c, x84, x85_c, x86, x88, x89_c, x90_c, x91, x93_c, x94_c, x95, x96, x98, x99_c);
and (w90, x0, x1_c, x2_c, x4_c, x6, x9_c, x11_c, x13_c, x14_c, x16_c, x21_c, x23, x24_c, x27_c, x29, x32, x33_c, x36, x37_c, x38_c, x39, x40, x41, x42, x44_c, x45_c, x46_c, x47, x48_c, x51_c, x52, x54, x55_c, x56_c, x58, x61, x62_c, x63, x65_c, x66, x67, x69_c, x70_c, x72_c, x74_c, x75, x77_c, x79, x80_c, x81, x82, x83_c, x84_c, x87, x88, x90, x91, x93, x94_c, x95, x97_c, x98);
and (w91, x4, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w92, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x71_c, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w93, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x41_c, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w94, x13_c, x38_c, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w95, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38_c, x83_c);
and (w96, x49, x85, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w97, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w98, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w99, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w100, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w101, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91, x92_c, x93_c, x95_c, x96, x98, x99);
and (w102, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x70_c, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w103, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w104, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w105, x4_c, x10, x15, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w106, x5, x10, x16, x21_c, x22, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w107, x0, x1, x2_c, x3, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w108, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78, x82, x83, x93_c, x97_c);
and (w109, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w110, x0, x3, x10, x13, x14, x15, x16_c, x22, x26, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w111, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80, x82, x83, x93_c, x97_c);
and (w112, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x90_c, x91, x96, x97_c, x98, x99);
and (w113, x0_c, x1, x2, x3, x4, x5_c, x6_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16, x17_c, x18, x19, x20_c, x21_c, x22_c, x23, x24, x25_c, x27, x28_c, x29, x30, x31, x32_c, x33, x35, x36_c, x37, x38_c, x39_c, x41, x42, x43, x44, x45, x46, x48, x49, x50_c, x51, x52, x53, x54, x55_c, x56, x57_c, x58, x59_c, x61_c, x62, x64_c, x65_c, x66_c, x67_c, x68, x70_c, x71, x72, x74, x75_c, x77_c, x78, x79_c, x81, x82, x83_c, x84, x85, x86, x87_c, x88, x91_c, x92_c, x93_c, x95, x96, x97_c, x98, x99);
and (w114, x0, x2_c, x3_c, x5_c, x7_c, x8, x9, x13_c, x16, x17_c, x20, x21, x23, x24, x25_c, x29_c, x32, x33_c, x34_c, x35, x39, x40_c, x41_c, x42, x44_c, x45, x46_c, x48_c, x49, x51_c, x52, x53, x55_c, x56, x58_c, x59_c, x60, x62, x65, x66, x67_c, x70, x71, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80_c, x86_c, x89, x93_c, x96, x99);
and (w115, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x57_c, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w116, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w117, x1, x2_c, x3_c, x8, x10_c, x11_c, x16_c, x17_c, x18_c, x19_c, x20, x21_c, x22, x23, x25, x27, x28, x29, x30_c, x31_c, x32_c, x33_c, x35, x36_c, x37_c, x42_c, x43_c, x45_c, x46, x50_c, x54_c, x55, x60_c, x62, x63_c, x64, x66_c, x68, x69_c, x72, x73, x75, x78_c, x84, x85_c, x89_c, x90, x94, x96_c, x99);
and (w118, x0_c, x4_c, x11, x14_c, x16, x17, x24_c, x25_c, x28, x29, x36_c, x37_c, x39_c, x51, x53, x55, x58, x59, x61, x69_c, x71_c, x74_c, x75, x76_c, x78_c, x79_c, x81, x82_c, x84, x87, x88, x95_c, x97_c, x98_c, x99);
and (w119, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x53_c, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w120, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x77, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w121, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w122, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90_c, x93_c, x97_c);
and (w123, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w124, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w125, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w126, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x84_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w127, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x69_c, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w128, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w129, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x39, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w130, x1, x2_c, x6, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w131, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w132, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w133, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x74_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w134, x13_c, x22, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w135, x0, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w136, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x34, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w137, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94, x95, x96, x97, x98);
and (w138, x0_c, x1_c, x3, x4, x7, x9_c, x12_c, x13_c, x16, x26, x27_c, x30, x32, x34_c, x35_c, x39, x43, x45_c, x48, x49_c, x50_c, x52, x55_c, x58, x59, x66, x67, x71, x74_c, x77, x83, x85_c, x88_c, x89, x90_c, x92, x95_c, x97);
and (w139, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w140, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x85_c, x86_c, x87, x88_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w141, x13_c, x14_c, x27_c, x40, x82, x90_c, x96, x98, x99_c);
and (w142, x2_c, x11, x16_c, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w143, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x50_c, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w144, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x51_c, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w145, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x91_c, x95, x96, x97, x99_c);
and (w146, x12_c, x32, x63_c, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w147, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9, x10, x11_c, x12_c, x13, x14, x15, x17_c, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28, x29_c, x30_c, x31_c, x32, x33_c, x36_c, x37_c, x38, x39_c, x40_c, x42_c, x43_c, x44, x45, x46_c, x47, x48_c, x49, x50, x51_c, x52, x53, x54, x55, x57_c, x58_c, x59, x60_c, x61, x62, x63, x64_c, x65, x66_c, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80, x81, x82_c, x83_c, x84_c, x85, x86, x87_c, x88, x89, x90, x91, x92, x93_c, x94, x95, x96, x98_c, x99_c);
and (w148, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w149, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w150, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86, x89, x93, x97_c, x98_c, x99_c);
and (w151, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w152, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x56_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w153, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w154, x0, x2, x3, x6_c, x10_c, x11, x12, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w155, x3_c, x5, x8, x15, x16_c, x19, x20_c, x21_c, x25_c, x26_c, x28, x31_c, x32, x33_c, x35_c, x36, x37, x44, x47_c, x48, x50, x56_c, x59_c, x64_c, x67, x68, x77_c, x80_c, x81, x86, x90, x91_c, x92, x94_c, x96, x98);
and (w156, x0_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w157, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x59_c, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w158, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w159, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x67, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w160, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w161, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w162, x0_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w163, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w164, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w165, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x23_c, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w166, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x80_c, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w167, x0, x2, x3_c, x4_c, x5, x6, x7, x8, x9_c, x10_c, x11, x12, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20, x21_c, x23, x24, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38_c, x39, x40, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47, x48, x49, x50_c, x51, x52_c, x53, x54, x55_c, x56_c, x57, x58, x59_c, x60, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68, x69, x70_c, x71, x72, x73_c, x74_c, x75, x76, x77_c, x78, x80, x81, x82_c, x83_c, x84_c, x85_c, x86, x87, x88_c, x90, x91_c, x92, x93, x94, x95, x96, x97, x98);
and (w168, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61_c, x83_c);
and (w169, x0_c, x1_c, x2_c, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w170, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w171, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w172, x12_c, x32, x48_c, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w173, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x73_c, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w174, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x37, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w175, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w176, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x44, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w177, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x37, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w178, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w179, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91, x92_c, x93, x97_c);
and (w180, x0, x1_c, x2, x3_c, x7, x8_c, x9_c, x10, x11, x12_c, x13, x14_c, x15_c, x17_c, x19_c, x20, x22, x23_c, x24_c, x25, x26, x27, x29_c, x30, x31_c, x32, x34, x35, x39, x40, x41, x42, x43, x44, x46_c, x47_c, x48, x49_c, x51, x52, x53_c, x54, x55_c, x56, x57_c, x58, x59_c, x60, x61_c, x62_c, x63, x64_c, x67_c, x68, x69, x70, x71, x72_c, x74_c, x75_c, x77_c, x78_c, x79, x80, x82, x83, x84_c, x85, x87, x88_c, x89, x91, x92, x94, x95_c, x96_c, x99_c);
and (w181, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w182, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74_c, x77_c, x80_c, x84_c, x90_c, x96, x98, x99_c);
and (w183, x3_c, x5, x6, x8, x16, x17_c, x21_c, x23_c, x26, x27, x34_c, x36, x38_c, x54, x57_c, x58_c, x61, x63, x66, x67, x69_c, x71_c, x73_c, x77, x79, x93_c, x95, x97_c, x98_c);
and (w184, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x23_c, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w185, x2_c, x3, x4_c, x6_c, x7_c, x8, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w186, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x67, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w187, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x31, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w188, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x35, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w189, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51_c, x83_c);
and (w190, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x72_c, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w191, x0_c, x1, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w192, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w193, x7_c, x8_c, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w194, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w195, x0_c, x1, x2, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w196, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x13_c, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w197, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w198, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x90_c, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w199, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w200, x13_c, x14_c, x37_c, x39_c, x45_c, x48_c, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w201, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82_c, x85, x89, x93, x97_c, x98_c, x99_c);
and (w202, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91, x93_c, x95_c, x96, x98, x99);
and (w203, x8, x21_c, x23, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w204, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x45, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w205, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w206, x5, x10, x16, x21_c, x31_c, x32, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w207, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w208, x0, x1_c, x2_c, x4, x6_c, x8_c, x13, x14_c, x17_c, x20, x23_c, x27, x28_c, x29, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x39_c, x46_c, x47_c, x48_c, x50, x51, x52, x53, x54, x55_c, x57, x59_c, x61_c, x62, x63_c, x64_c, x66, x68, x69, x70_c, x71, x73_c, x74, x75, x77_c, x78_c, x79, x80_c, x83, x84_c, x87, x92_c, x93, x94_c, x95, x99);
and (w209, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x90_c, x93_c, x96_c, x97_c, x98, x99);
and (w210, x1_c, x17, x19_c, x30_c, x42_c, x43, x44_c, x55, x56, x59, x64_c, x66_c, x73, x82_c, x86_c, x90_c);
and (w211, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x29, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w212, x0_c, x1, x2_c, x3_c, x4, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x21, x22, x23_c, x24, x26, x27_c, x28, x29, x30_c, x31, x32, x33, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x43_c, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51, x52, x53, x54_c, x55_c, x56, x58_c, x59_c, x60_c, x61, x62_c, x63, x64, x65_c, x66, x67_c, x68, x69, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79_c, x81_c, x82, x83_c, x84_c, x85_c, x86, x87, x88, x89, x90_c, x91_c, x92, x93_c, x94, x95_c, x96, x97_c, x98_c, x99);
and (w213, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w214, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94, x95, x96_c, x97, x98, x99);
and (w215, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w216, x1_c, x2, x4, x5_c, x6_c, x9_c, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w217, x2_c, x3_c, x5, x7, x8, x9_c, x10_c, x12, x13, x16, x17, x20_c, x22_c, x24_c, x26_c, x27_c, x28, x29_c, x30_c, x31_c, x32, x33_c, x35_c, x36, x41_c, x42, x43, x44, x45_c, x46, x47, x50, x51, x52, x53, x57_c, x58_c, x60_c, x62_c, x63, x64, x65, x66, x69_c, x72_c, x73, x76, x78, x80, x81_c, x83, x85_c, x87, x89_c, x95, x98_c, x99_c);
and (w218, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x37_c, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w219, x3, x5_c, x18, x21_c, x33_c, x39_c, x76, x77_c, x94);
and (w220, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w221, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w222, x12_c, x32, x40_c, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w223, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x81, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w224, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x91_c, x92, x95, x97_c);
and (w225, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w226, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13_c, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w227, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w228, x5_c, x9, x27, x61_c, x76, x80, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w229, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w230, x0_c, x1, x3_c, x4_c, x5, x6_c, x7_c, x10_c, x11, x12_c, x13, x14_c, x15_c, x16, x17_c, x18_c, x19, x21_c, x23_c, x24, x27, x28_c, x29, x30, x32_c, x34_c, x35, x36_c, x37, x38, x39, x40, x41_c, x42, x43_c, x44, x45, x46, x47_c, x48, x50, x51, x52, x54, x55, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x65, x66, x67_c, x69_c, x70, x71_c, x72_c, x73_c, x75, x76_c, x78, x80_c, x81, x82, x83, x84, x85, x86, x87_c, x88, x89_c, x90_c, x91, x92_c, x93, x94, x95_c, x96, x97_c, x99);
and (w231, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x50, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w232, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w233, x0, x1_c, x3, x5_c, x6, x7_c, x8_c, x10, x11, x12_c, x13, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30_c, x31_c, x32, x33, x36_c, x39, x40, x41, x42, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x52_c, x53, x54, x55_c, x57_c, x58_c, x59, x60, x61_c, x63, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71, x72, x73_c, x74_c, x75, x77_c, x78_c, x79, x80_c, x82, x83, x84, x85_c, x87_c, x88, x89_c, x90_c, x91, x92_c, x93, x94_c, x96_c, x97, x98, x99);
and (w234, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x80_c, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w235, x3_c, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w236, x1_c, x3, x10, x12, x16, x26_c, x29, x30, x42, x44, x47, x53_c, x54, x57_c, x59_c, x61_c, x68, x69, x74, x81_c, x87, x91);
and (w237, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92, x96_c, x97_c, x98, x99_c);
and (w238, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x95, x96, x97_c, x98, x99_c);
and (w239, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w240, x12_c, x32, x84, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w241, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x59, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w242, x49, x73, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w243, x12_c, x32, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w244, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w245, x12_c, x40, x56, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w246, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87_c, x95, x99);
and (w247, x0, x1, x2_c, x7, x10, x12_c, x14_c, x20, x21_c, x23_c, x24_c, x25, x26, x29, x33, x36, x37, x38, x41, x49, x54_c, x62_c, x72, x74, x76_c, x77, x80, x81_c, x83, x86_c, x87, x89_c, x94_c, x95, x96, x97, x98);
and (w248, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w249, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x21, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w250, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x84, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w251, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w252, x13_c, x14_c, x37_c, x39_c, x45_c, x50_c, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w253, x0_c, x5, x20, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w254, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w255, x13_c, x49_c, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w256, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x80, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w257, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60_c, x83_c);
and (w258, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x41, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w259, x0, x1_c, x2_c, x3, x4, x5_c, x10, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w260, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w261, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w262, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w263, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w264, x3_c, x4, x5_c, x8, x9_c, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w265, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x54_c, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w266, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86_c, x95, x99);
and (w267, x0, x2, x3, x6_c, x10_c, x11, x13_c, x17_c, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w268, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x21, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w269, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w270, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w271, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97, x99);
and (w272, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91, x92, x93_c, x94, x95_c, x96, x98, x99);
and (w273, x0, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w274, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54_c, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w275, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w276, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23_c, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w277, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w278, x0_c, x1_c, x2_c, x5_c, x6_c, x7, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18, x19_c, x20, x21_c, x22_c, x23_c, x24_c, x25, x26, x27_c, x28_c, x29_c, x31_c, x33, x34_c, x35, x36_c, x37_c, x39, x41_c, x45_c, x46, x48, x49_c, x50_c, x52_c, x53_c, x54, x55_c, x56_c, x57, x59_c, x60_c, x63_c, x64, x66, x67, x70_c, x71_c, x72, x73, x74_c, x75, x76, x77, x78, x79, x81_c, x82_c, x83_c, x84_c, x86, x88, x90_c, x92_c, x93, x94, x96_c, x97_c, x98);
and (w279, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91, x92, x94_c, x95, x96_c, x98, x99_c);
and (w280, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x80_c, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w281, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x72_c, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w282, x0_c, x2_c, x3, x5_c, x6, x7, x8, x9, x10, x11_c, x14, x15_c, x16, x17, x20, x21, x22, x23_c, x25, x26, x27, x28, x29, x30_c, x32, x33, x34, x36, x38_c, x40_c, x42_c, x43_c, x44, x46_c, x47, x48_c, x49_c, x50_c, x51_c, x52, x53, x54, x55, x60_c, x61, x62_c, x63_c, x64, x65, x67, x68_c, x72_c, x73, x74_c, x77, x78_c, x79, x80, x84_c, x85, x86, x88, x90_c, x92, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w283, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w284, x0, x1_c, x2, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w285, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w286, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w287, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w288, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x90_c, x91, x95, x96, x98, x99);
and (w289, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w290, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w291, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w292, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x82_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w293, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x90_c, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w294, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x50_c, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w295, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x25_c, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w296, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79, x82, x83, x93_c, x97_c);
and (w297, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88, x90, x91_c, x95, x96, x97, x99_c);
and (w298, x3_c, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w299, x0, x2, x4_c, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w300, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x61_c, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w301, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x58_c, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w302, x35, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w303, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w304, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w305, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w306, x0_c, x1_c, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10, x11, x12_c, x13_c, x14_c, x15, x16, x17, x18, x19_c, x20, x21_c, x22_c, x23, x24, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31, x32_c, x33, x34, x35_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x43_c, x44, x46, x47, x48, x49, x50_c, x51, x53_c, x54, x55_c, x56_c, x57, x58_c, x59, x60_c, x61_c, x62, x63_c, x64_c, x66, x67, x68, x69_c, x70, x71, x72, x73_c, x74_c, x75, x76, x77, x78, x79_c, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88_c, x89_c, x90, x91, x92, x93, x94_c, x95, x96, x97_c, x98_c);
and (w307, x2_c, x11, x29_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w308, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w309, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w310, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85, x90_c, x93_c, x95_c, x96, x98, x99);
and (w311, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x39, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w312, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
assign w313 = x94;
and (w314, x0_c, x2_c, x4, x6, x8_c, x11_c, x13_c, x16_c, x17_c, x18_c, x19, x21_c, x22_c, x23, x24_c, x28, x29, x32_c, x33_c, x34, x35, x36, x37, x38_c, x39, x40, x41_c, x43, x45, x46_c, x47, x48, x49, x50, x51_c, x53_c, x55_c, x56_c, x59_c, x60_c, x61, x62, x64, x65, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x73, x75, x76_c, x77, x78_c, x81, x82, x83_c, x84_c, x85, x87, x89, x90_c, x91, x92, x93, x94_c, x95_c, x96_c, x97, x98, x99);
and (w315, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w316, x0, x2, x3, x6_c, x10_c, x11, x13_c, x14_c, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w317, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w318, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w319, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w320, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x61_c, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w321, x12_c, x32, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w322, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w323, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w324, x4_c, x5_c, x7_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w325, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x77_c, x90_c, x93_c, x97_c);
and (w326, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w327, x0, x1_c, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w328, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x47, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w329, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w330, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x14, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w331, x5, x7_c, x15_c, x17, x31, x34, x38_c, x40, x41, x47, x67, x69_c, x70_c, x76, x79_c, x85_c, x87_c, x88_c, x91, x94);
and (w332, x0, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15, x17_c, x18, x19, x20_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x34, x35, x36, x37_c, x38_c, x39, x40, x41_c, x43, x44_c, x45_c, x46, x47, x48, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57_c, x58_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x66, x67, x68_c, x69_c, x70, x71, x72, x73_c, x74_c, x75_c, x76, x77, x78, x79_c, x80_c, x81_c, x82, x83, x84, x85_c, x86_c, x87, x88, x89_c, x90, x91, x92_c, x93, x94, x95, x96, x97, x98_c, x99_c);
and (w333, x3_c, x8_c, x12, x14_c, x15_c, x18, x19, x21, x22, x23, x24, x25, x28, x31, x32, x34, x37_c, x41_c, x43_c, x44_c, x46, x50, x51, x52, x53, x54_c, x55_c, x56, x57, x62_c, x63, x64, x68, x71_c, x73_c, x78_c, x79, x80, x81_c, x85_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w334, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x65, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w335, x6, x17_c, x20_c, x21_c, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w336, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x93, x94_c, x95, x96_c, x98, x99_c);
and (w337, x0, x2, x7_c, x8_c, x11, x13_c, x18, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w338, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x60, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w339, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w340, x13_c, x14_c, x37_c, x39_c, x43, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w341, x8, x21_c, x25_c, x27_c, x34, x36, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w342, x0_c, x2_c, x3, x6_c, x10_c, x11, x13_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w343, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w344, x12_c, x16, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w345, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x59_c, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w346, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w347, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w348, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x94, x95_c, x97_c);
and (w349, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w350, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w351, x0_c, x1, x2, x5_c, x7, x8_c, x9_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w352, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w353, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w354, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w355, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63_c, x83_c);
and (w356, x12_c, x32, x91, x96_c, x97_c, x98, x99);
and (w357, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73_c, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w358, x1, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w359, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x80, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w360, x5_c, x9, x27, x61_c, x71_c, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w361, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w362, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w363, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x84, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w364, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w365, x2_c, x11, x29_c, x41, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w366, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x87_c, x89_c, x90, x93, x94_c, x96, x97);
and (w367, x12_c, x40, x78, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w368, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92_c, x97_c);
and (w369, x0_c, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w370, x0, x1_c, x3, x5_c, x7, x10, x26_c, x27_c, x31, x33_c, x34_c, x39_c, x44_c, x50_c, x52, x53, x54_c, x57, x58, x65_c, x90_c, x92_c, x95_c, x96, x97);
and (w371, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w372, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72, x75_c, x77, x82, x83, x93_c, x97_c);
and (w373, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w374, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57_c, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w375, x4_c, x5_c, x7_c, x8, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w376, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x18, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w377, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57_c, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w378, x1, x2_c, x4_c, x6, x7_c, x8_c, x11, x14_c, x17, x18_c, x20, x21_c, x22, x23, x24, x25_c, x26, x27_c, x29_c, x30_c, x32, x35_c, x37, x38_c, x42_c, x44_c, x45_c, x47_c, x48_c, x50, x52, x53_c, x54, x56, x57_c, x58_c, x62_c, x63, x65, x66_c, x67, x68_c, x69, x70_c, x72_c, x74, x77_c, x78_c, x79, x80_c, x82_c, x85, x86_c, x87_c, x88, x89_c, x90, x91, x92_c, x95_c, x96);
and (w379, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x32, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w380, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w381, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w382, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x81_c, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w383, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x37, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w384, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85_c, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w385, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w386, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w387, x6, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w388, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67, x75_c, x77, x82, x83, x93_c, x97_c);
and (w389, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w390, x26_c, x58_c, x62_c, x70, x94);
and (w391, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x30, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w392, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w393, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w394, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w395, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60_c, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w396, x1_c, x2, x7, x13, x19_c, x20_c, x23_c, x24_c, x29_c, x35, x39_c, x45_c, x54, x61_c, x69, x70_c, x71_c, x73_c, x79, x81, x85_c, x90, x92, x97, x99_c);
and (w397, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78, x85, x89, x93, x97_c);
and (w398, x1, x3_c, x5, x10_c, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w399, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x94, x95, x96, x97_c, x98_c, x99_c);
and (w400, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w401, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41, x82, x90_c, x96, x98, x99_c);
and (w402, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x59_c, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w403, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w404, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x82, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w405, x0_c, x1_c, x2, x3, x4, x5, x6_c, x7_c, x8, x9, x10_c, x12, x13, x14, x15, x16_c, x17_c, x18_c, x19, x20, x21, x22, x23, x24, x26_c, x27_c, x29, x30_c, x31_c, x32_c, x33, x34_c, x35, x36_c, x37, x38_c, x39_c, x40, x41, x42, x43, x44, x45, x46, x47, x48_c, x50, x51_c, x52_c, x53, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61, x62, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73_c, x74, x75, x76, x77, x78, x79_c, x80, x81, x82_c, x84_c, x85_c, x86_c, x87, x88_c, x89, x90, x91_c, x92_c, x93, x94, x95, x96_c, x98_c, x99_c);
and (w406, x2_c, x4_c, x5, x9, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w407, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91, x92, x93_c, x94, x95_c, x98, x99_c);
and (w408, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w409, x33_c, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w410, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w411, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w412, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x64_c, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w413, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x34_c, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w414, x5, x10, x16, x21_c, x34_c, x35, x38, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w415, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x95_c, x97_c);
and (w416, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92, x93_c, x95_c, x96, x97, x98_c, x99_c);
and (w417, x34, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w418, x1, x5_c, x16, x17, x19_c, x26_c, x30_c, x35_c, x37, x39, x40_c, x46, x48_c, x49_c, x52, x63_c, x72, x73, x74_c, x76_c, x79, x81_c, x83_c, x84_c, x89_c);
and (w419, x0_c, x1_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w420, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w421, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51_c, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w422, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65_c, x83_c);
and (w423, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w424, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x89_c, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w425, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w426, x73, x78, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w427, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x16, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w428, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x58_c, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w429, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80, x82, x83, x93_c, x97_c);
and (w430, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w431, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w432, x8, x30_c, x38, x41_c, x49, x56_c, x87, x92_c);
and (w433, x3, x5, x7, x12_c, x21_c, x25, x28, x35, x39, x41, x47, x48, x56, x57_c, x59, x65_c, x68_c, x71, x76_c, x79_c, x81, x88_c, x89, x90_c, x95_c, x97_c, x98, x99_c);
and (w434, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x91_c, x93, x95_c, x96_c, x99);
and (w435, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w436, x4_c, x5_c, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w437, x0, x1, x2_c, x4, x5_c, x6, x7_c, x8, x9, x10, x11, x13, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x30, x31_c, x32, x33_c, x34, x35, x36_c, x37, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46, x47_c, x48, x49_c, x50_c, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62_c, x63_c, x64, x65_c, x66, x67_c, x68_c, x69_c, x70, x71, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x79, x80, x81_c, x82, x83_c, x84, x86, x87, x88, x89, x90_c, x91, x92, x93, x94_c, x95, x96, x97, x98_c, x99);
and (w438, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w439, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w440, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x32, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w441, x0_c, x1_c, x2, x3_c, x5_c, x6, x7, x9_c, x10, x11_c, x12_c, x13_c, x15, x16, x17_c, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25_c, x26_c, x27, x28, x29, x30_c, x31, x32, x33, x34_c, x35_c, x36_c, x37, x39_c, x40, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54_c, x55_c, x56, x57, x58_c, x59, x60, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70_c, x71_c, x72, x73, x74, x75, x76, x77_c, x78, x79_c, x81_c, x83_c, x85_c, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98, x99_c);
and (w442, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w443, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w444, x2_c, x3_c, x4_c, x6_c, x9, x10_c, x12_c, x13, x14, x15_c, x17_c, x18_c, x19_c, x21_c, x24_c, x25, x26, x27, x29_c, x30, x32_c, x33, x35, x36, x37_c, x39, x40_c, x45_c, x48_c, x50_c, x52_c, x56, x58, x59, x60_c, x61, x65_c, x67_c, x68_c, x69_c, x70, x71, x72, x73, x77_c, x78_c, x79, x81_c, x83_c, x85, x88_c, x89, x90, x91_c, x92_c, x93, x95_c, x97_c);
and (w445, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x66, x75_c, x77, x82, x83, x93_c, x97_c);
and (w446, x9_c, x17_c, x26, x27, x28_c, x31_c, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w447, x13_c, x14_c, x37_c, x39_c, x45_c, x47_c, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w448, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x96, x98, x99);
and (w449, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w450, x0_c, x1_c, x3_c, x5_c, x7_c, x10, x11_c, x14, x19_c, x21, x23, x24_c, x29, x30, x31, x34, x36, x39_c, x40, x41, x44_c, x46_c, x47, x49_c, x50_c, x59, x63_c, x66, x68_c, x70_c, x73_c, x75_c, x77_c, x78, x79, x80_c, x81, x83_c, x84, x86_c, x88, x90_c, x93_c, x94_c, x96, x97, x98);
and (w451, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x13, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w452, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91, x92, x93_c, x97_c);
and (w453, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x82, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w454, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x29_c, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w455, x0, x1_c, x4_c, x5_c, x6_c, x7_c, x8, x9_c, x10, x11, x13, x15, x16_c, x17, x19, x20_c, x21, x22, x23, x24, x25, x27_c, x28, x29, x30, x31_c, x33, x34, x35, x36_c, x39, x41_c, x43, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50_c, x51, x52_c, x53, x55, x56, x57, x58, x60, x61_c, x63, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x72, x73_c, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81, x82, x83, x84, x85_c, x86_c, x89_c, x91_c, x92_c, x93, x94_c, x95, x96_c);
and (w456, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91, x92_c, x94_c, x97_c);
and (w457, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w458, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x89_c, x91_c, x92, x93, x94, x95_c, x97_c);
and (w459, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x72_c, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w460, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x57_c, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w461, x1_c, x7_c, x8_c, x9_c, x13_c, x15_c, x17, x19, x20, x24, x25, x28, x31, x43_c, x44_c, x48, x49, x53, x54_c, x55_c, x60_c, x61, x62, x63_c, x64_c, x68_c, x72, x76_c, x79_c, x82, x85_c, x88, x89_c, x96_c);
and (w462, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w463, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92_c, x93_c, x95_c, x96, x98, x99);
and (w464, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w465, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x49, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w466, x1, x2, x3, x4, x5, x6, x7, x8_c, x9_c, x10, x12, x13, x14_c, x15, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24, x25_c, x26_c, x28_c, x29_c, x30, x31, x32, x33, x36, x39, x40_c, x41_c, x42_c, x43_c, x44, x45, x46, x47, x49_c, x51, x52_c, x53, x54, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66_c, x67, x68, x69, x70, x71, x72_c, x73, x76_c, x77_c, x78_c, x79, x80_c, x82_c, x84, x85_c, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94, x95, x96, x97, x98_c, x99);
and (w467, x0, x3, x10, x13, x14, x15, x16_c, x22, x33, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w468, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x92_c, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w469, x0, x3, x10, x13, x14, x15, x16_c, x22, x32, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w470, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w471, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29_c, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w472, x0, x12_c, x40, x82, x90_c, x96, x98, x99_c);
and (w473, x0_c, x1, x2, x3_c, x4, x5, x6, x7, x8_c, x9, x10_c, x11, x12, x13, x14, x16_c, x18_c, x19_c, x20, x21_c, x22_c, x23, x24_c, x25, x26_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34, x36_c, x37, x38, x40, x41_c, x42, x44_c, x45_c, x46_c, x47_c, x48, x49_c, x50, x51_c, x54_c, x55, x56_c, x58_c, x60_c, x61_c, x63_c, x65_c, x66, x68, x70_c, x71, x72, x74_c, x76_c, x77, x79, x81_c, x82_c, x83, x84, x85, x86_c, x88_c, x90, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w474, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w475, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14_c, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w476, x5_c, x9, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w477, x0, x1, x2, x3_c, x4, x5, x6_c, x7_c, x8_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x24, x25_c, x26, x27_c, x28, x29, x30, x31, x32_c, x33, x34, x35_c, x36, x37, x38, x39, x40, x41_c, x42_c, x43, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56, x57, x58, x59_c, x60_c, x61_c, x62, x63_c, x64, x65_c, x66, x67, x68, x69, x70_c, x71_c, x72, x73, x74, x75, x76_c, x77_c, x78_c, x79, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x88, x89_c, x90, x91, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w478, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w479, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w480, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w481, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94, x95, x96_c, x97_c, x98, x99_c);
and (w482, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w483, x5, x10, x16, x21_c, x27, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w484, x0_c, x1, x2_c, x3_c, x4, x5, x6_c, x7, x8, x9, x10_c, x11_c, x12_c, x13, x14_c, x15_c, x16, x17_c, x18_c, x19, x20, x21_c, x22_c, x23_c, x24, x25, x26_c, x27, x28_c, x30_c, x31, x32_c, x33_c, x34_c, x36_c, x37_c, x39_c, x40, x41_c, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50_c, x51, x52_c, x53, x54, x55_c, x56_c, x57_c, x58, x60, x61, x62_c, x63, x64, x65_c, x66, x67, x68_c, x69, x70, x71_c, x72, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84, x85_c, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94_c, x95_c, x96_c, x97, x98, x99_c);
and (w485, x1_c, x7, x8, x12, x15, x17, x20_c, x23, x24_c, x27_c, x32_c, x35_c, x36_c, x39, x40_c, x43, x49, x51_c, x53, x55_c, x59_c, x63_c, x65, x69_c, x70, x72, x76_c, x82_c, x83_c, x85_c, x87, x89_c, x92, x93, x96_c, x97);
and (w486, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w487, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w488, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w489, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w490, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x36_c, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w491, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x77, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w492, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92_c, x93_c, x97_c);
and (w493, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80_c, x81, x84, x85, x95, x99);
and (w494, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w495, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x56, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w496, x13_c, x49, x53_c, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w497, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15_c, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w498, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w499, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w500, x1_c, x2_c, x3, x4, x5, x11_c, x13, x14_c, x17, x18_c, x23, x24_c, x25_c, x27, x28, x31_c, x32_c, x33_c, x34_c, x38, x40, x42, x43_c, x44_c, x45, x48_c, x51, x52, x53_c, x54, x56, x57_c, x59_c, x62, x66, x67, x69, x73, x81, x82_c, x87, x90_c, x91_c, x92, x94_c, x97, x98, x99);
and (w501, x4_c, x10, x15_c, x19, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w502, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w503, x1, x2, x5_c, x7, x12_c, x16_c, x19, x26, x30, x31, x32_c, x36, x38_c, x40_c, x42_c, x43_c, x48_c, x49_c, x56_c, x60_c, x62_c, x65_c, x70_c, x73_c, x75_c, x79, x81_c, x84_c, x85, x87_c, x88, x91_c, x93_c, x94, x98_c);
and (w504, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78_c, x82, x83, x93_c, x97_c);
and (w505, x0, x2_c, x3_c, x4_c, x5_c, x6, x7, x9, x12_c, x14, x16, x17, x18, x19, x20_c, x21, x26_c, x28_c, x29, x35, x38, x41, x42_c, x43_c, x46_c, x47, x48, x51, x52, x53, x54_c, x55_c, x56, x58, x59_c, x60_c, x63_c, x64_c, x65, x66_c, x68_c, x71, x72, x73_c, x74_c, x77, x78_c, x79_c, x81_c, x83_c, x86, x90_c, x91, x93, x95, x97, x98);
and (w506, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w507, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x93_c, x94_c, x95, x96_c, x98, x99_c);
and (w508, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x55_c, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w509, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w510, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x91_c, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w511, x8, x21_c, x25_c, x27_c, x32_c, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w512, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x58, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w513, x0_c, x1, x2, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w514, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w515, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w516, x65_c, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w517, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x83_c, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w518, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x44, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w519, x2_c, x8_c, x9_c, x32, x33_c, x37_c, x39_c, x40, x54_c, x56_c, x57, x68_c, x70, x75, x79, x87, x89, x91_c, x94, x97);
and (w520, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w521, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w522, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w523, x12_c, x32, x58_c, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w524, x0_c, x5, x7, x12_c, x13, x14, x16_c, x19, x20, x24, x27, x29_c, x31, x33_c, x36, x37, x38, x40, x41_c, x42_c, x43, x44_c, x45_c, x47_c, x50_c, x53, x65, x67_c, x68, x69_c, x70, x71, x75, x78_c, x79_c, x81_c, x82, x83_c, x84_c, x86_c, x92, x93_c, x94, x95, x96_c, x98);
and (w525, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x65, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w526, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w527, x8, x21_c, x25_c, x27_c, x31_c, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w528, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14_c, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w529, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22_c, x40, x82, x90_c, x96, x98, x99_c);
and (w530, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x84, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w531, x0_c, x2_c, x6_c, x7, x8_c, x10, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w532, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w533, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w534, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w535, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x53_c, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w536, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x55, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w537, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w538, x4_c, x10, x13_c, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w539, x1_c, x3, x5, x6, x9, x13, x19_c, x20_c, x28_c, x31_c, x32_c, x35, x40, x41, x43_c, x46, x48, x51_c, x55_c, x56, x57_c, x61_c, x63, x64, x65_c, x66, x67, x68, x70, x71_c, x72_c, x73_c, x74, x77_c, x87_c, x89, x90, x91_c, x97_c, x98, x99_c);
and (w540, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84_c, x90_c, x93_c, x97_c);
and (w541, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74_c, x81, x84, x85, x95, x99);
and (w542, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w543, x0, x2, x3_c, x4, x6_c, x7_c, x10, x11_c, x18, x19, x20_c, x21, x24, x25_c, x26_c, x27_c, x28, x30_c, x32_c, x33, x35_c, x37, x39, x40_c, x42_c, x43_c, x46_c, x47_c, x48, x49, x52, x54_c, x55, x56_c, x58_c, x59, x61_c, x62_c, x63, x67_c, x69_c, x70_c, x72, x73, x74_c, x75_c, x77, x78_c, x79, x80_c, x81, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x92_c, x94_c, x95_c, x96_c, x97_c);
and (w544, x0, x2_c, x3_c, x5, x6, x8, x10_c, x11_c, x13_c, x14, x15, x17_c, x18, x20_c, x23, x24, x25, x27, x28_c, x29, x31_c, x34_c, x35_c, x36, x38_c, x39, x43, x45_c, x48, x49_c, x51_c, x52_c, x54_c, x55, x56_c, x57_c, x60, x61, x62, x63, x65_c, x67, x70, x71_c, x72_c, x73, x74, x76_c, x78, x82, x85, x88, x90, x91_c, x92_c, x93_c, x96_c, x97, x98_c, x99);
and (w545, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x28_c, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w546, x0_c, x1_c, x3_c, x5_c, x6_c, x7_c, x9_c, x10, x12, x13, x14_c, x15_c, x16, x17, x18_c, x20_c, x21, x23_c, x24, x25_c, x29, x31, x32, x33_c, x34, x35_c, x36_c, x38, x41_c, x42, x44_c, x45, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x54_c, x55_c, x56_c, x60, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x70_c, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x79, x81_c, x82_c, x84, x85_c, x87_c, x88, x89, x90_c, x92_c, x93_c, x94_c, x95_c, x97, x98_c);
and (w547, x49, x87, x88, x92, x94_c, x95_c, x96, x97_c);
and (w548, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w549, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w550, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w551, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91);
and (w552, x1, x3, x5, x6_c, x7_c, x9_c, x12, x16_c, x20, x21_c, x22, x24_c, x28_c, x29, x34_c, x42_c, x45, x46_c, x54_c, x57_c, x58_c, x63, x69, x70, x73, x78_c, x83, x84_c, x88_c, x89, x96_c, x98_c, x99_c);
and (w553, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w554, x0, x3, x10, x13, x14, x15, x16_c, x20_c, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w555, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x66, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w556, x0, x1_c, x4_c, x9, x10_c, x12_c, x13_c, x15_c, x16_c, x19_c, x20, x21, x22, x23, x28, x29_c, x31_c, x32_c, x34_c, x35_c, x37_c, x38, x44, x47, x50, x53_c, x55, x56, x57, x61, x62_c, x64, x65_c, x66_c, x69, x70, x74_c, x77_c, x78, x80_c, x82, x85, x87, x90_c, x93, x94_c, x96_c, x97_c, x98);
and (w557, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x75, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w558, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w559, x3_c, x5, x6_c, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w560, x8, x13_c, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w561, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w562, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w563, x0_c, x3, x5_c, x10_c, x14_c, x19, x25, x26_c, x29, x30_c, x33_c, x37, x39_c, x42_c, x43, x44_c, x49_c, x51, x61, x64_c, x67_c, x68, x69_c, x72, x78_c, x92_c, x97_c, x99);
and (w564, x12_c, x32, x72_c, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w565, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x46, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w566, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x13, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w567, x5_c, x9, x27, x50_c, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w568, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x29, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w569, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x87, x90, x91_c, x95, x96, x97, x99_c);
and (w570, x4_c, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w571, x3_c, x4, x5, x8, x9_c, x10_c, x12_c, x17, x18_c, x19, x20_c, x21, x22, x23_c, x24, x26, x28, x29_c, x30, x31, x35, x37, x42_c, x45_c, x47_c, x48, x50_c, x51_c, x53, x55, x56, x57_c, x58_c, x59, x61, x62, x63, x65_c, x66_c, x67_c, x69, x73_c, x74_c, x75_c, x76, x79, x82_c, x85_c, x86_c, x89, x93);
and (w572, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x41_c, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w573, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x79, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w574, x0_c, x1, x2, x3, x4, x5_c, x6, x7_c, x8, x9, x10, x11_c, x12, x14, x16_c, x17, x18, x19, x20, x21, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29_c, x30, x31, x32, x33, x34_c, x36_c, x37, x38_c, x39, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48_c, x49, x50_c, x51_c, x52_c, x53, x54, x55, x56, x57_c, x59, x60, x62_c, x63, x64_c, x65, x66, x67_c, x68, x69, x70_c, x71, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x79_c, x80_c, x81, x82, x83, x84, x85, x86_c, x87, x88, x89_c, x90, x91, x92, x93, x94, x95, x96_c, x97, x98_c, x99_c);
and (w575, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w576, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w577, x0, x1_c, x13, x22, x24, x25_c, x30, x43, x46_c, x48, x54_c, x60_c, x61_c, x65, x66, x67_c, x75_c, x81_c, x83, x87_c, x89, x98, x99_c);
and (w578, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x57_c, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w579, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x82, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w580, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91, x92, x93_c, x94, x96, x97);
and (w581, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w582, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w583, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x53_c, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w584, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w585, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x86, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w586, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x74_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w587, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x92, x95_c, x97_c);
and (w588, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w589, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w590, x1, x2_c, x6_c, x15, x16, x47, x57, x79_c, x95_c, x97);
and (w591, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x93_c, x95_c, x96, x97_c, x98, x99_c);
and (w592, x4, x5, x6_c, x7, x8_c, x9_c, x10, x12_c, x13_c, x14_c, x15_c, x16, x17, x18, x19, x20_c, x21, x22_c, x23_c, x24, x26_c, x27_c, x28, x29, x30, x31_c, x32, x33_c, x34, x35_c, x36, x38, x39_c, x40, x41_c, x42_c, x43_c, x45, x46, x48_c, x49_c, x50, x52, x53, x54, x55_c, x57, x58, x59_c, x60_c, x61_c, x62, x63_c, x64, x66, x67, x68_c, x69, x71, x74_c, x75_c, x76, x77_c, x78_c, x81_c, x82_c, x83, x84_c, x85_c, x86_c, x87_c, x88, x89, x90_c, x92, x94, x95_c, x96, x97_c, x98_c, x99);
and (w593, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w594, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w595, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62_c, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w596, x5, x10, x16, x17_c, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w597, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w598, x6_c, x7_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w599, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w600, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55_c, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w601, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x57_c, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w602, x0, x1, x2, x3, x4, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13, x14_c, x16, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26_c, x27, x28_c, x29, x30, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48_c, x49_c, x50, x51_c, x52, x53, x54_c, x55_c, x56, x57_c, x58, x59_c, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80, x81_c, x82_c, x83, x84_c, x85, x86, x87_c, x88, x89, x90, x91_c, x92_c, x94_c, x95, x96_c, x97, x98, x99);
and (w603, x8, x21_c, x22, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w604, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w605, x0_c, x1, x2, x3_c, x4, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w606, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x61, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w607, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77_c, x79, x90_c, x93_c, x97_c);
and (w608, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w609, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w610, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w611, x0, x1_c, x2, x3_c, x4, x5_c, x6, x8, x9, x11, x12_c, x13_c, x15_c, x16, x17, x19, x20_c, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x40_c, x41, x42, x43, x44_c, x45_c, x47, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56_c, x57, x58, x59, x60, x61_c, x62, x63, x64, x65, x68, x69, x70, x71_c, x72, x73, x75_c, x77, x79_c, x80_c, x81, x82_c, x83_c, x85_c, x86_c, x87_c, x88_c, x89_c, x92, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w612, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69_c, x83_c);
and (w613, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w614, x6, x17_c, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w615, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w616, x11, x12_c, x15, x17_c, x18, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w617, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x40_c, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w618, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w619, x0_c, x1, x2, x3_c, x5, x6, x7_c, x8, x9_c, x10_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28_c, x29_c, x30, x31_c, x32, x34, x35_c, x37, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45, x46_c, x47, x49, x50_c, x51_c, x52_c, x53_c, x54, x56, x58_c, x59_c, x61, x62_c, x63, x64, x65, x66, x67, x68_c, x69, x70_c, x71, x72_c, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84, x85, x86, x87_c, x88, x89, x90, x91, x92_c, x95, x96, x97_c, x98, x99_c);
and (w620, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88, x90_c, x93_c, x95_c, x96, x97_c, x98, x99);
and (w621, x2_c, x3_c, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w622, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x86, x88_c, x90_c, x91, x92, x95, x97_c);
and (w623, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w624, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w625, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w626, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w627, x49, x58_c, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w628, x3, x13, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w629, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w630, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x18, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w631, x3, x5_c, x14, x38_c, x39_c, x42_c, x45_c, x51_c, x54, x64_c);
and (w632, x3_c, x4, x5_c, x7, x25_c, x36, x38, x46_c, x49, x51_c, x54, x61, x63_c, x76_c, x77_c, x78, x89, x91, x93);
and (w633, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90);
and (w634, x0, x1_c, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w635, x0, x2_c, x3_c, x5, x7_c, x9, x10_c, x11, x12, x13_c, x15, x18, x20_c, x23_c, x25, x26, x28, x31, x33_c, x37, x39, x40_c, x42, x47, x48, x49, x51, x52_c, x53, x54_c, x55_c, x57_c, x60, x62_c, x64, x67, x75, x76_c, x78, x80, x81_c, x82, x84_c, x86, x87_c, x88, x90, x95_c, x97, x98);
and (w636, x5_c, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w637, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w638, x4, x5_c, x9_c, x26_c, x35_c, x37, x42, x45, x49, x80, x84);
and (w639, x4_c, x10, x15_c, x22_c, x24_c, x27, x30_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w640, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91, x92_c, x94, x96, x99);
and (w641, x6, x16, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w642, x0_c, x4_c, x7, x8_c, x12, x13_c, x14_c, x18_c, x19_c, x21, x37_c, x38, x46_c, x47, x48, x49_c, x52_c, x53, x55_c, x57, x58_c, x61, x63, x66_c, x67, x68_c, x72, x75_c, x83, x84, x86, x87_c, x89, x91, x97_c);
and (w643, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w644, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93, x96, x98, x99_c);
and (w645, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w646, x2, x3_c, x9, x13, x14, x15, x20, x35, x37, x38_c, x39_c, x40_c, x41_c, x43_c, x44_c, x45_c, x46_c, x47_c, x51, x53, x55, x57_c, x59, x61, x64_c, x65, x66_c, x72_c, x76_c, x82_c, x84_c, x85, x86, x88_c, x92_c, x93);
and (w647, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w648, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w649, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x62, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w650, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23_c, x40, x82, x90_c, x96, x98, x99_c);
and (w651, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x55_c, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w652, x0, x4_c, x15_c, x19_c, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w653, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w654, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w655, x47_c, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w656, x9_c, x17_c, x19_c, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w657, x0, x1, x2_c, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12, x13_c, x14, x15, x16_c, x17_c, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x28, x29, x30_c, x31_c, x32, x33_c, x34_c, x35_c, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x45, x46, x47_c, x48, x49_c, x50, x51_c, x52_c, x53, x54, x55_c, x56, x57, x58_c, x59_c, x60_c, x61, x62, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73, x74, x75_c, x76_c, x77, x78_c, x79_c, x81_c, x82_c, x83, x85_c, x86, x87, x88, x89_c, x90, x91, x92_c, x93, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w658, x0, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w659, x2_c, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w660, x0_c, x1_c, x2, x3, x4, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x14, x15_c, x16_c, x17_c, x19_c, x20, x21, x22_c, x23, x24_c, x25, x26, x27, x29, x30_c, x31, x32_c, x33, x34, x35_c, x36_c, x38, x39, x40_c, x41_c, x42, x43, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x54, x55_c, x57_c, x58, x59_c, x60_c, x61_c, x62, x63_c, x64_c, x65, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74, x76_c, x77, x78_c, x79_c, x80, x81, x82_c, x83_c, x84, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95_c, x97_c, x98, x99);
and (w661, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w662, x8, x21_c, x25_c, x27_c, x31_c, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w663, x3, x13, x16, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w664, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w665, x0, x1, x2, x4, x8, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w666, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x26_c, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w667, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w668, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30_c, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w669, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w670, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81, x82, x83, x93_c, x97_c);
and (w671, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x72_c, x81, x84, x85, x95, x99);
and (w672, x5_c, x9, x20, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w673, x1_c, x24_c, x31_c, x39_c, x47, x55_c, x58, x63_c, x73_c, x78_c, x80_c, x85, x89_c, x92_c, x94);
and (w674, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x88_c, x89, x91, x93_c, x94_c, x95_c, x96, x97, x98);
and (w675, x0, x1_c, x2_c, x3_c, x4_c, x5, x6_c, x7, x8_c, x9, x10_c, x11_c, x12, x13, x14_c, x15_c, x16, x17_c, x18_c, x19, x20, x21_c, x22_c, x23_c, x24, x25, x26, x27_c, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34_c, x35, x36_c, x37, x38, x39, x40, x41_c, x42_c, x43, x44_c, x45_c, x46_c, x47, x49, x50_c, x51, x52_c, x54, x56_c, x57_c, x58_c, x59, x60_c, x61, x62, x63_c, x65, x66_c, x67_c, x68, x69_c, x70, x71, x72, x73_c, x74, x75_c, x76_c, x77, x78, x79_c, x81, x82_c, x83, x84_c, x85_c, x86, x87_c, x88_c, x90, x91, x92_c, x93_c, x94, x95, x96, x97, x98, x99_c);
and (w676, x0_c, x1_c, x2, x3_c, x4_c, x6, x7, x8, x9, x10_c, x12_c, x14_c, x15_c, x16, x17_c, x19_c, x20, x23, x24, x25, x27, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x37_c, x38_c, x39, x40_c, x41, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x51, x52_c, x54, x56, x57, x58, x60, x61_c, x62, x63, x67, x69, x72_c, x73, x77, x78, x79_c, x80, x81_c, x83, x84_c, x85, x87_c, x88, x90, x92_c, x93, x94, x95, x97_c, x98_c);
and (w677, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x28, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w678, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w679, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w680, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x41_c, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w681, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w682, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x81, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w683, x5_c, x9, x27, x33_c, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w684, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w685, x12_c, x31, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w686, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w687, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w688, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x23, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w689, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81_c, x83_c);
and (w690, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x63, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w691, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x32_c, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w692, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w693, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w694, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w695, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w696, x0_c, x3_c, x4_c, x6, x7_c, x8, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w697, x49, x51_c, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w698, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w699, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x71_c, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w700, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x67_c, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w701, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w702, x0, x3_c, x13_c, x15, x16_c, x17, x19_c, x23_c, x25, x46_c, x50_c, x54_c, x58_c, x59, x67_c, x72_c, x76_c, x85, x86, x94, x99_c);
and (w703, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x69_c, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w704, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x40_c, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w705, x0_c, x3_c, x4_c, x6, x7_c, x10_c, x12_c, x40, x82, x90_c, x96, x98, x99_c);
and (w706, x1_c, x8_c, x19_c, x20, x29_c, x36_c, x51, x52, x54_c, x55_c, x63, x66_c, x68, x74_c, x84, x86_c, x88_c, x94_c);
and (w707, x1_c, x16, x32_c, x49, x64, x80);
and (w708, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72_c, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w709, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w710, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w711, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x17_c, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w712, x0_c, x1_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w713, x1, x3_c, x5, x9_c, x10_c, x13, x15_c, x17, x18, x19, x21_c, x22, x24_c, x25_c, x26, x27_c, x29_c, x30_c, x31_c, x32_c, x33, x39, x41_c, x42, x43_c, x44_c, x46, x47_c, x49, x50, x51_c, x53, x54, x55, x57, x58_c, x60, x61_c, x62_c, x65, x66, x67, x68_c, x69, x70_c, x71_c, x73_c, x75_c, x76, x77_c, x80, x81, x82_c, x86_c, x87_c, x88_c, x90_c, x91_c, x93_c, x95_c, x97_c, x98_c, x99);
and (w714, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90_c, x93_c, x95_c, x96, x98, x99);
and (w715, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x18_c, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w716, x31_c, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w717, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w718, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w719, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w720, x49, x88_c, x92, x94_c, x95_c, x96, x97_c);
and (w721, x10_c, x11, x13, x15, x17, x20, x27_c, x31_c, x44, x46, x55_c, x68, x78_c, x81, x88_c, x91_c, x93_c);
and (w722, x5, x10, x16, x20, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w723, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x33_c, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w724, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w725, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w726, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w727, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w728, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76, x79, x90_c, x93_c, x97_c);
and (w729, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x55, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w730, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w731, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97);
and (w732, x3, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w733, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w734, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x22_c, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w735, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99);
and (w736, x1, x2_c, x3_c, x5_c, x6_c, x7, x10_c, x12_c, x13_c, x14_c, x15, x16_c, x17, x21_c, x22_c, x25, x26, x27_c, x32_c, x34_c, x36, x38, x40_c, x41_c, x42, x43, x45, x46_c, x48_c, x49, x50, x51_c, x52, x53, x55, x57, x58, x61_c, x62, x64_c, x65_c, x66, x67_c, x68_c, x69_c, x70, x76_c, x77, x78, x79_c, x80, x81, x82_c, x84, x85_c, x87, x88_c, x89_c, x93, x94, x96_c, x99_c);
and (w737, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w738, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w739, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x90, x93_c, x97_c);
and (w740, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x43, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w741, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w742, x0, x2, x5_c, x6_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w743, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x15, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w744, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w745, x1, x4_c, x5_c, x6, x7, x8, x10_c, x11_c, x12, x14_c, x15_c, x17_c, x18, x19_c, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x31, x32, x33, x36, x37_c, x38_c, x39_c, x40, x41_c, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x52_c, x54, x55, x56, x57_c, x58, x59_c, x60, x61_c, x62_c, x63_c, x64, x66, x67, x68, x69, x72_c, x73_c, x74_c, x76, x78, x79_c, x81_c, x83_c, x84, x85, x86_c, x87, x88, x89, x90, x91_c, x93, x94, x95_c, x96_c, x97_c);
and (w746, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w747, x0, x3, x10, x13, x14_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w748, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w749, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22_c, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w750, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w751, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w752, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x27_c, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w753, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x89_c, x93, x97_c);
and (w754, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w755, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x35, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w756, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x52, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w757, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x12, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w758, x0_c, x1, x3_c, x6_c, x7, x8, x10, x12, x13_c, x14, x15, x16, x18, x20_c, x21, x23_c, x24_c, x25, x26, x29_c, x35_c, x37, x39, x41_c, x42_c, x43_c, x44, x45, x48_c, x49, x50, x51, x52_c, x54_c, x55, x56, x57, x59, x61, x62_c, x64, x65, x66, x68_c, x70, x71, x72_c, x75_c, x77, x78, x79, x80, x81, x85_c, x87, x88, x89, x90_c, x91, x93_c, x96, x98_c, x99);
and (w759, x0_c, x3, x5, x7, x9, x11_c, x12, x13, x14_c, x16_c, x18_c, x19, x20, x21_c, x22_c, x24_c, x25, x26, x28, x32_c, x34, x35_c, x39_c, x40, x44, x45_c, x46, x47, x48, x49, x50, x51_c, x54, x57, x58_c, x62, x64_c, x65_c, x68, x70_c, x73_c, x76, x77_c, x79, x83_c, x84_c, x85, x87, x89_c, x91, x92_c, x93, x94_c, x96, x97_c, x98, x99_c);
and (w760, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x69_c, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w761, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x64, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w762, x12_c, x40, x82, x90_c, x99);
and (w763, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w764, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w765, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x47_c, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w766, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x41, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w767, x0_c, x2, x3_c, x6, x7, x8_c, x11_c, x12, x14, x15_c, x17, x22, x25_c, x26_c, x27, x32_c, x39_c, x42, x48_c, x50, x56_c, x64_c, x65_c, x67_c, x78, x80, x83, x84_c, x85_c, x86, x89, x90_c, x92_c, x94_c);
and (w768, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x9, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w769, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w770, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w771, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x21, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w772, x12_c, x32, x79, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w773, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x48, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w774, x0, x1_c, x2_c, x3, x5_c, x6_c, x7_c, x8_c, x11, x12_c, x13, x17_c, x19_c, x20, x23_c, x24_c, x25_c, x26, x28, x30, x31, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x41, x42, x43, x44, x45_c, x46, x47_c, x48, x49_c, x52_c, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61_c, x62, x64, x65_c, x68_c, x70_c, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80_c, x82_c, x83, x84, x85, x87_c, x88_c, x89, x90, x91_c, x93_c, x94, x95, x96_c, x97_c, x99_c);
and (w775, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w776, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w777, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w778, x0_c, x1_c, x2, x3_c, x4, x5, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14_c, x15, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30_c, x31_c, x32, x33, x34_c, x35, x37_c, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47_c, x48_c, x49_c, x50, x51, x52, x53_c, x55_c, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64, x65_c, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92_c, x93, x94, x95, x96, x97_c, x98_c, x99);
and (w779, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w780, x0, x1_c, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w781, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28_c, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w782, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81, x84_c, x85_c, x97_c);
and (w783, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x15, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w784, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
assign w785 = x20_c;
and (w786, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14, x15_c, x16, x17_c, x18, x19_c, x20, x21_c, x22, x23, x24, x25_c, x26, x27, x28_c, x29, x30, x31_c, x32, x33_c, x34_c, x35, x36_c, x37_c, x38_c, x39_c, x40, x41, x42_c, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56, x57, x58, x59_c, x60_c, x61_c, x62, x63, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x81, x82_c, x83, x84, x85, x86_c, x87, x88_c, x89, x90_c, x91, x92, x93, x94, x95, x96_c, x97_c, x98, x99);
and (w787, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x61, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w788, x0_c, x3_c, x7, x9, x11, x17, x21_c, x24, x32_c, x36_c, x38, x43, x44, x45_c, x47_c, x53, x58_c, x61, x62, x65_c, x69, x73, x81_c, x84_c, x87_c, x91_c, x92);
and (w789, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w790, x42, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w791, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x23_c, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w792, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w793, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x27_c, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w794, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w795, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w796, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68, x72_c, x81, x84, x85, x95, x99);
and (w797, x5, x10, x16, x21_c, x34_c, x35_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w798, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w799, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w800, x12_c, x14, x20_c, x26, x44, x53_c, x74, x99);
and (w801, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w802, x49, x82_c, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w803, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46, x73_c, x76, x85, x89, x93, x97_c);
and (w804, x6, x9, x11, x15, x16_c, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w805, x5_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w806, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w807, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w808, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x45_c, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w809, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x54_c, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w810, x0, x1_c, x2, x4_c, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w811, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w812, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92, x93_c, x97_c);
and (w813, x28_c, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w814, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91_c, x92, x93, x94_c, x95_c, x97_c);
and (w815, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w816, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w817, x0, x1, x3, x6, x7_c, x9, x10, x11_c, x12_c, x13, x14_c, x15_c, x16_c, x17_c, x18, x19, x21_c, x23, x24_c, x25, x26, x27_c, x28, x30_c, x32, x33, x34_c, x36_c, x37, x40, x41_c, x43, x44, x45_c, x46, x47, x49_c, x51_c, x53, x54, x55, x56, x57, x59_c, x60_c, x62, x63_c, x65, x67_c, x68, x70_c, x71, x73, x75_c, x76, x77, x79, x81_c, x82, x83_c, x85, x86, x87, x88, x89_c, x91, x92, x94, x96, x98, x99_c);
and (w818, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x87, x88, x91, x93_c);
and (w819, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76_c, x83_c);
and (w820, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w821, x0_c, x3_c, x4_c, x6, x7_c, x10, x11_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w822, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x24, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w823, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x47, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w824, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w825, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w826, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w827, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w828, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w829, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x58_c, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w830, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x69_c, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w831, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w832, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w833, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x90_c, x91, x96, x97, x98_c, x99_c);
and (w834, x0_c, x2_c, x3, x4_c, x5_c, x6, x7, x11_c, x13_c, x19_c, x20_c, x21_c, x22, x24, x27_c, x28_c, x29_c, x30, x32_c, x33, x34, x35_c, x36, x37_c, x38, x39, x40, x41_c, x42, x44_c, x46_c, x52_c, x54_c, x55, x57, x60, x62_c, x63, x65, x68_c, x69, x70_c, x71_c, x72_c, x73, x75, x78, x79, x80_c, x81_c, x83, x84, x86_c, x88_c, x89_c, x91, x92_c, x93_c, x95, x96, x97);
and (w835, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w836, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80, x90_c, x93_c, x97_c);
and (w837, x72, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w838, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x93, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w839, x0_c, x1_c, x3, x4_c, x5, x6_c, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w840, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x62_c, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w841, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x64_c, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w842, x0_c, x2_c, x4_c, x7_c, x9, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w843, x8, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w844, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69, x75_c, x77, x82, x83, x93_c, x97_c);
and (w845, x0, x2, x5_c, x6, x7, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w846, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x96, x97_c, x98, x99_c);
and (w847, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w848, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x93, x94_c, x95, x96_c, x98, x99_c);
and (w849, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w850, x0, x3, x10, x13_c, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w851, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x81_c, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w852, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x82, x83, x93_c, x97_c);
and (w853, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w854, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w855, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w856, x0_c, x1, x2, x3_c, x5, x6_c, x7_c, x8, x10_c, x11_c, x12, x13, x14, x15_c, x16_c, x17, x18, x19, x20, x21_c, x22, x23, x25_c, x28_c, x29, x30_c, x31_c, x32_c, x33, x34, x36_c, x37, x38, x39_c, x40, x41, x42, x43_c, x44_c, x45_c, x46, x48, x49_c, x51, x53, x54_c, x55_c, x56, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x66, x67_c, x68, x69, x70, x71_c, x72_c, x74_c, x77, x78_c, x79_c, x80, x81, x82_c, x83, x84_c, x85, x86, x87, x88_c, x89_c, x90, x91_c, x93, x95_c, x96, x97, x98_c);
and (w857, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w858, x2, x6, x7_c, x9_c, x10_c, x11, x14, x18, x22_c, x23, x24_c, x28_c, x29, x30, x31, x34_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x41_c, x43_c, x44_c, x47_c, x48, x49, x50_c, x51, x53, x55_c, x56_c, x58_c, x59, x62, x63_c, x64_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x75, x77_c, x80, x81_c, x82_c, x83_c, x84_c, x85, x87, x89_c, x90, x91, x93, x96, x97_c, x98_c);
and (w859, x1, x2_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w860, x0, x1_c, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w861, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x89_c, x90_c, x92_c, x93, x95_c);
and (w862, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87_c, x90_c, x93_c, x97_c);
and (w863, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w864, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w865, x34, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w866, x0, x4_c, x15_c, x21_c, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w867, x2, x3, x8, x11, x12_c, x18, x22_c, x24, x40, x47_c, x50_c, x55, x60, x65_c, x70_c, x78, x81_c, x85_c, x86_c, x97_c);
and (w868, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x92_c, x93, x94_c, x95, x96_c, x98, x99_c);
and (w869, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w870, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w871, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w872, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x41_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w873, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x97);
and (w874, x0_c, x1, x2, x3_c, x4, x5_c, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w875, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x66_c, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w876, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w877, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x70_c, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w878, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67, x71_c);
and (w879, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w880, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x60_c, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w881, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81, x82, x83, x93_c, x97_c);
and (w882, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w883, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13_c, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w884, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w885, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x42_c, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w886, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91_c, x93_c, x95_c, x96, x98, x99);
and (w887, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x32_c, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w888, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x50_c, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w889, x0, x1, x2_c, x3_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w890, x2, x6_c, x43_c);
and (w891, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x86, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w892, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50_c, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w893, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w894, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w895, x3, x5_c, x8, x14_c, x15, x30_c, x35, x36, x38, x39, x40, x49, x61, x62_c, x76_c);
and (w896, x0, x1, x2, x4, x7, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w897, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w898, x9, x13, x17, x19, x28_c, x37, x42, x47_c, x54, x64_c, x85, x86, x89_c, x91_c, x93_c, x96);
and (w899, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w900, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x87, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w901, x7, x9_c, x11_c, x40_c, x49, x54_c, x59, x66, x72, x74, x84_c, x86, x90, x92_c, x99_c);
and (w902, x0_c, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w903, x8, x12_c, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w904, x0, x1, x2, x3_c, x4, x5, x6_c, x7, x8_c, x9, x12, x13, x15, x16, x18_c, x19_c, x20, x22, x23_c, x24, x26_c, x27_c, x28_c, x29_c, x30, x32, x34, x35_c, x36_c, x37, x38_c, x40, x42, x43, x44, x45_c, x46_c, x47_c, x48, x50_c, x51_c, x56, x57_c, x59_c, x60_c, x61, x62, x63_c, x64, x66_c, x67, x70_c, x72, x74_c, x75, x77, x78, x80_c, x81, x82, x83, x86, x88, x89_c, x91, x92, x93, x94_c, x95, x96_c, x97_c, x99_c);
and (w905, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w906, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x42, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w907, x4_c, x9_c, x14, x16_c, x25_c, x34_c, x55_c, x61, x75_c, x76, x83_c, x86_c, x88, x89_c);
and (w908, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w909, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x94, x95, x96_c, x97, x98, x99_c);
and (w910, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x54, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w911, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x32, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w912, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w913, x13, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w914, x2, x4_c, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w915, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x81_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w916, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x75_c, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w917, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x65, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w918, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w919, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w920, x12_c, x40, x82, x90_c, x93_c, x94_c, x95, x96_c, x98, x99_c);
and (w921, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w922, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w923, x9_c, x16, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w924, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w925, x25_c, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w926, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x9, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w927, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x80, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w928, x66_c, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w929, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x87_c, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w930, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42_c, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w931, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w932, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66_c, x75, x84_c, x85_c, x97_c);
and (w933, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w934, x49, x72, x73, x79, x90_c, x93_c, x97_c);
and (w935, x13_c, x49, x64, x71, x72_c, x79, x87_c, x90, x93_c, x97_c);
and (w936, x6, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w937, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x84, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w938, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x35, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w939, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41_c, x83_c);
and (w940, x23, x62, x66_c, x67, x70_c);
and (w941, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w942, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w943, x8, x21_c, x25_c, x26_c, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w944, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x90, x91, x92, x95, x97_c);
and (w945, x3_c, x7_c, x12, x13_c, x14, x16, x18, x19_c, x23, x24_c, x25, x29, x34_c, x37, x38, x40, x43_c, x45, x48_c, x50_c, x52_c, x57, x59_c, x61_c, x64_c, x66, x68, x69_c, x74, x82, x84_c, x87_c, x89, x90_c, x92, x94_c, x97_c);
and (w946, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w947, x12_c, x40, x81_c, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w948, x0_c, x3_c, x4_c, x6, x7_c, x10, x11_c, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w949, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62, x73_c, x76, x85, x89, x93, x97_c);
and (w950, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w951, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w952, x0, x1, x2_c, x6_c, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w953, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w954, x2, x3, x5_c, x6_c, x10, x11, x12_c, x13, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x23_c, x24_c, x26, x28, x31_c, x32, x33_c, x34, x38, x39_c, x41_c, x43, x44_c, x45_c, x46_c, x47, x51_c, x52, x54, x62_c, x65, x66_c, x67_c, x68, x71, x73_c, x75_c, x77, x79, x80_c, x81, x82, x84, x85_c, x86_c, x87_c, x89_c, x90, x91, x92, x94, x96, x97_c, x98_c);
and (w955, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24_c, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w956, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w957, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w958, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c, x98, x99_c);
and (w959, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x22, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w960, x12_c, x33_c, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w961, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x61, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w962, x3, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w963, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69, x75_c, x77, x82, x83, x93_c, x97_c);
and (w964, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22_c, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w965, x10, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w966, x0_c, x1_c, x3_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w967, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x43, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w968, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w969, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w970, x3_c, x7_c, x9_c, x12_c, x15, x17, x18_c, x22, x24_c, x27_c, x30, x32, x33_c, x34_c, x35_c, x37_c, x39_c, x40_c, x41_c, x45_c, x46_c, x47, x49, x52_c, x54_c, x55, x56_c, x58, x59_c, x60_c, x61, x62, x64_c, x66, x68, x72_c, x73, x74_c, x76, x77, x80, x81, x86_c, x88, x90, x92, x95_c, x96);
and (w971, x5, x10, x16, x21_c, x32_c, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w972, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w973, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x74, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w974, x1, x2_c, x5_c, x6_c, x9_c, x14_c, x17, x18_c, x19, x24, x27_c, x31, x37_c, x40, x41, x46, x49, x51, x61, x68, x90_c, x96_c);
and (w975, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w976, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x33_c, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w977, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w978, x3, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w979, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w980, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w981, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w982, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w983, x6, x17_c, x20_c, x24_c, x25_c, x26, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w984, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w985, x1_c, x4_c, x7_c, x9, x10, x13_c, x14_c, x15_c, x16, x17_c, x20, x25_c, x28_c, x29, x30_c, x31_c, x32_c, x34, x35_c, x36_c, x37_c, x39, x43, x47, x49_c, x52_c, x53_c, x54_c, x56, x65_c, x66, x68_c, x70_c, x73_c, x74, x78_c, x80, x84, x89, x90, x93_c, x99);
and (w986, x2_c, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w987, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w988, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x19, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w989, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87, x93_c, x97_c);
and (w990, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w991, x0_c, x1_c, x3_c, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w992, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x32, x83_c);
and (w993, x0, x1, x2_c, x8, x9_c, x10, x17, x21, x26_c, x27_c, x29_c, x34_c, x40, x41_c, x42_c, x45_c, x48, x49, x50, x54_c, x56, x59, x62, x65_c, x66, x68_c, x75_c, x78_c, x80_c, x82, x85_c, x89_c, x92, x93, x94, x95, x96, x97, x98, x99_c);
and (w994, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w995, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w996, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x13_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w997, x5_c, x9, x27, x61_c, x76, x88_c, x97);
and (w998, x1, x3, x4_c, x5, x7, x8_c, x10_c, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w999, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88_c, x89, x93, x97_c);
and (w1000, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8_c, x10, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1001, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x86, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1002, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x65_c, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1003, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1004, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1005, x13_c, x49, x54, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w1006, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x80_c, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1007, x2_c, x5_c, x7, x8_c, x12, x15_c, x16, x18_c, x21, x22_c, x23_c, x24, x26_c, x30, x33, x38_c, x40, x45_c, x47_c, x54_c, x55, x56, x57_c, x60, x63_c, x64, x65, x67, x68_c, x69_c, x70_c, x75_c, x78_c, x79, x80_c, x83_c, x87, x88_c, x90, x92_c, x98);
and (w1008, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1009, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1010, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1011, x3_c, x4, x7, x9_c, x23, x25, x26_c, x28_c, x30, x44_c, x49, x50_c, x52, x53, x54, x57_c, x61_c, x65_c, x68, x70, x73, x78, x80_c, x81, x82_c, x83, x89, x90_c, x92, x93_c, x95, x96_c);
and (w1012, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x91, x93_c, x95_c, x96, x98, x99);
and (w1013, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x41, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1014, x2, x5_c, x9, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1015, x15, x17_c, x25_c, x27, x32_c, x33_c, x34, x38, x40_c, x42_c, x43_c, x44_c, x66_c, x68, x74_c, x75, x89_c, x97_c);
and (w1016, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1017, x4, x42_c, x63_c);
and (w1018, x8, x19, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1019, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1020, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x57, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1021, x2, x4_c, x5, x6, x7_c, x9_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1022, x2, x4_c, x7, x9, x10, x13, x14, x15, x16, x17_c, x18_c, x19_c, x20, x24_c, x26, x27, x29, x30, x32_c, x35, x36, x37, x40_c, x41, x43_c, x46_c, x48, x50_c, x52_c, x53_c, x55, x56_c, x60_c, x62, x66_c, x67_c, x69, x73, x75, x76, x77, x78_c, x79, x82, x83, x84_c, x85, x86, x87, x89_c, x91, x92_c, x93_c, x94_c, x97_c, x99);
and (w1023, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1024, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x28_c, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1025, x9_c, x17_c, x26, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1026, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1027, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1028, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x45_c, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1029, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1030, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1031, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x77, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1032, x0_c, x1, x2_c, x3, x4_c, x5, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1033, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x41_c, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1034, x6, x11_c, x15, x16_c, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w1035, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1036, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42_c, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1037, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x69, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1038, x0_c, x1_c, x3, x5, x6_c, x7_c, x8_c, x9, x10, x11_c, x12_c, x13_c, x14_c, x19_c, x21, x22, x23, x26_c, x27_c, x28, x29, x30, x31, x33_c, x34, x35, x36_c, x38_c, x39_c, x40, x41_c, x44_c, x45_c, x48, x49, x51, x52, x54_c, x55_c, x56_c, x57_c, x58_c, x60_c, x62, x63_c, x64_c, x66, x67_c, x69, x70, x72, x73_c, x74_c, x76, x77_c, x79, x82, x89_c, x90_c, x91, x92, x94_c, x96_c, x98);
and (w1039, x1_c, x2_c, x11, x12_c, x15, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1040, x2_c, x11, x29_c, x68, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1041, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37, x71_c);
and (w1042, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1043, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x30_c, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1044, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1045, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1046, x0_c, x2, x7, x9, x14, x22, x26, x28_c, x40, x54, x58, x59_c, x60, x62_c, x65_c, x70, x84_c, x98);
and (w1047, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79, x80_c, x82, x83_c, x84);
and (w1048, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88, x89_c, x90, x91_c, x92_c, x93, x94, x95, x96_c, x98, x99_c);
and (w1049, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1050, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x45_c, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1051, x2_c, x11, x29_c, x90, x93_c, x95_c, x96, x98, x99);
and (w1052, x11, x12_c, x15, x17_c, x23_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1053, x49, x72, x73_c, x74, x75, x76_c, x77_c, x79, x90_c, x93_c, x97_c);
and (w1054, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29, x40, x82, x90_c, x96, x98, x99_c);
and (w1055, x4, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1056, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1057, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1058, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90_c, x95, x99);
and (w1059, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x45, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1060, x0_c, x1_c, x2_c, x3_c, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14, x15, x17, x18_c, x19, x20_c, x21_c, x22, x23, x24, x25, x26_c, x27_c, x28_c, x29_c, x30_c, x31, x32, x33_c, x34_c, x35, x36, x37, x38, x39_c, x40_c, x41_c, x42, x43, x44_c, x45_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55, x56_c, x58_c, x59, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69, x70_c, x71, x72_c, x73, x74, x75, x76_c, x77_c, x78, x79_c, x80_c, x81, x82, x83_c, x84, x85, x86, x87, x89, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97, x98_c, x99);
and (w1061, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91_c, x93_c, x95_c, x96, x98, x99);
and (w1062, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x25, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1063, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90, x93_c, x97_c);
and (w1064, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1065, x9_c, x17_c, x18_c, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1066, x4, x6, x8, x11, x15_c, x16_c, x17, x20, x23, x25_c, x26_c, x29_c, x34_c, x36, x38_c, x41, x47_c, x49_c, x53, x55_c, x64, x67_c, x70_c, x75, x78, x85, x88, x90_c, x91, x92, x95_c);
and (w1067, x0, x5_c, x10, x12, x18_c, x23, x24_c, x25_c, x27, x36, x37_c, x44, x49_c, x53_c, x64_c, x65, x78, x82, x87_c, x93, x95, x97_c, x98);
and (w1068, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x56, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1069, x8, x21_c, x25_c, x27_c, x34, x39_c, x41_c, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1070, x0, x1, x2_c, x3, x4, x6_c, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1071, x2_c, x3_c, x4, x6, x7, x8, x10, x11, x14, x16, x17, x19, x21, x25, x27, x28, x30_c, x31, x32_c, x35_c, x36_c, x37_c, x39, x40, x42, x43_c, x44, x45, x46_c, x49, x50, x52_c, x54, x57, x58_c, x59, x60, x62, x65, x66, x68_c, x69_c, x72_c, x73_c, x82, x83, x84_c, x88_c, x89, x91_c, x92, x93, x97, x98);
and (w1072, x53, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1073, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1074, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x82, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1075, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x92_c, x93_c, x94, x95, x96_c, x97_c);
and (w1076, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x11_c, x12, x13, x15_c, x16_c, x17_c, x18, x19, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x27_c, x29, x30, x31, x32, x34_c, x36, x37_c, x38_c, x41, x42_c, x43_c, x44, x46, x49_c, x51, x53, x55, x56_c, x57, x58, x59_c, x60, x61_c, x64, x65, x66_c, x67_c, x70, x71, x72_c, x73_c, x74, x75, x76_c, x77, x78_c, x79, x80, x82_c, x83_c, x84_c, x85_c, x86, x87, x88, x89, x90, x92, x96_c, x97);
and (w1077, x73, x77, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1078, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x95_c, x96_c, x97, x98, x99_c);
and (w1079, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1080, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1081, x2_c, x3, x7, x11, x14, x16_c, x18_c, x19_c, x25, x38, x47_c, x48_c, x54_c, x55, x59, x60_c, x61_c, x67, x68, x69_c, x71_c, x72_c, x73, x75, x76_c, x79_c, x80, x84, x85_c, x87, x89_c, x90_c, x91, x93, x94, x95, x96_c, x98_c);
and (w1082, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1083, x68, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1084, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1085, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1086, x7, x9, x15, x17, x21_c, x24_c, x29, x34, x37_c, x42_c, x46, x50_c, x51, x55_c, x63, x64, x66, x67, x68, x69, x72_c, x73, x79_c, x83_c, x89, x92_c, x93, x97_c, x98, x99);
and (w1087, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20_c, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1088, x0, x3_c, x4_c, x5_c, x6, x7_c, x8_c, x11, x12_c, x13_c, x17, x20, x21, x22, x23, x24_c, x25_c, x27_c, x28_c, x29_c, x30, x31, x32_c, x35_c, x41, x42, x43_c, x45_c, x46, x47_c, x48, x52, x54_c, x55_c, x56_c, x58, x59, x62_c, x63, x64_c, x65, x66_c, x67, x69_c, x70, x71_c, x72, x76, x77_c, x78_c, x79_c, x80_c, x84, x87_c, x91_c, x92_c, x93_c, x95, x96_c, x98_c, x99);
and (w1089, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w1090, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56, x82, x90_c, x96, x98, x99_c);
and (w1091, x0_c, x3_c, x6, x11_c, x14, x15, x20, x22, x24, x25, x27_c, x29_c, x30_c, x33_c, x35, x39_c, x41_c, x44, x45_c, x46, x48_c, x51_c, x53, x55, x58_c, x60_c, x62_c, x63, x64, x65, x66_c, x67, x70_c, x72, x75_c, x85_c, x88, x89_c, x90, x91_c);
and (w1092, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1093, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1094, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x98_c, x99);
and (w1095, x0_c, x1, x2, x3_c, x4_c, x5_c, x7, x8_c, x9_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1096, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w1097, x0, x2, x3, x6_c, x8_c, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1098, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1099, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x73, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1100, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1101, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1102, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x59, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1103, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71_c, x83_c);
and (w1104, x0_c, x2_c, x4_c, x5, x7_c, x11_c, x12, x16_c, x17, x18, x19_c, x24, x25, x33_c, x35_c, x38, x40_c, x41_c, x42_c, x46_c, x47, x48, x50, x51, x56, x57_c, x65, x67_c, x68, x76_c, x81, x87_c, x88_c, x89, x95);
and (w1105, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1106, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x84_c, x85_c, x90, x96, x98, x99_c);
and (w1107, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1108, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1109, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1110, x2, x3, x7_c, x14_c, x17_c, x22, x23, x24, x26, x27, x31, x33, x35_c, x38, x39_c, x41, x42_c, x46, x48_c, x49, x54_c, x56, x57, x58_c, x62_c, x65_c, x71, x72, x79, x82_c, x84_c, x89_c, x90_c, x91_c, x97);
and (w1111, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x64_c, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1112, x12_c, x40, x76_c, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1113, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1114, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31_c, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1115, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x50, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1116, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1117, x13_c, x30_c, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w1118, x26, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1119, x8, x14_c, x16_c, x18, x22, x23_c, x27_c, x37, x38_c, x40, x51_c, x57, x62, x65_c, x70, x71_c, x72_c, x73_c, x76, x79_c, x83, x90);
and (w1120, x0_c, x1_c, x2_c, x3_c, x4_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13_c, x14, x15_c, x16, x17, x18, x19_c, x21_c, x22, x23, x25_c, x27, x28, x29_c, x30, x31, x32_c, x33, x34, x35, x36, x37_c, x38_c, x39, x41, x43, x44_c, x45_c, x46, x47, x48_c, x49, x51, x53, x54_c, x56_c, x58, x59, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69, x70, x71_c, x72_c, x73_c, x74_c, x75, x77, x78_c, x79, x81_c, x82_c, x83, x84_c, x85_c, x87_c, x89_c, x90, x91_c, x92_c, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w1121, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1122, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x65_c, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1123, x12_c, x40, x41_c, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1124, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1125, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x22_c, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1126, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x83_c);
and (w1127, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87_c, x88, x89_c, x90_c, x91_c, x92, x93_c, x95, x97_c);
and (w1128, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x42, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1129, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x91, x92_c, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w1130, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1131, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x64, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1132, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x13_c, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1133, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x50_c, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1134, x12_c, x40, x47, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1135, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1136, x17, x30, x38, x41_c, x72, x83_c, x91);
and (w1137, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1138, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1139, x0_c, x3, x12_c, x40, x82, x90_c, x96, x98, x99_c);
and (w1140, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1141, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x83_c);
and (w1142, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92_c);
and (w1143, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1144, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x85_c, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1145, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1146, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1147, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x64_c, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1148, x13_c, x14_c, x37_c, x39_c, x40, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1149, x0, x5_c, x6_c, x8, x9_c, x11_c, x12_c, x13, x21_c, x22, x24, x26_c, x28_c, x30, x35, x37_c, x40_c, x41_c, x42, x47_c, x48, x50, x51_c, x53, x55, x56_c, x60, x63, x64_c, x69_c, x80_c, x83, x84_c, x86_c, x88_c, x97_c);
and (w1150, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x48_c, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1151, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x80_c, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1152, x12_c, x40, x77, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1153, x37, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1154, x12_c, x14, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1155, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94_c);
and (w1156, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1157, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89, x91_c, x92);
and (w1158, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84_c, x93_c, x97_c);
and (w1159, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1160, x0_c, x1, x2, x3_c, x4, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1161, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1162, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1163, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x73, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1164, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1165, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1166, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1167, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57, x82, x90_c, x96, x98, x99_c);
and (w1168, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92_c, x94_c, x95_c, x97, x98, x99);
and (w1169, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x37, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1170, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1171, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x45, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1172, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x37, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1173, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1174, x0, x1_c, x2, x7_c, x8_c, x10_c, x13_c, x14, x15_c, x16_c, x17_c, x20_c, x21_c, x24, x25_c, x26_c, x28, x30_c, x32, x34, x38_c, x42_c, x43, x50, x53_c, x55, x57_c, x58_c, x59, x61_c, x62_c, x63_c, x64_c, x65, x67, x69_c, x70_c, x72_c, x73_c, x74_c, x77_c, x79_c, x87_c, x92, x94_c, x95_c, x96_c, x97);
and (w1175, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1176, x4_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w1177, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1178, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w1179, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1180, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1181, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x40, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1182, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x52_c, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1183, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x70_c, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1184, x0_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1185, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1186, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x75, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w1187, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1188, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1189, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78_c, x81, x84, x85, x95, x99);
and (w1190, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1191, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1192, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1193, x1_c, x2, x5_c, x6, x11_c, x12, x14, x15, x19_c, x26_c, x27, x30, x32_c, x35, x39, x41_c, x42_c, x43, x49, x55, x62_c, x63, x64_c, x67_c, x70_c, x71_c, x72, x75, x76, x79, x80_c, x82, x84, x85_c, x89, x90_c, x93, x96);
and (w1194, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1195, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x88_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1196, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1197, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1198, x6, x12, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1199, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1200, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x24, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1201, x0, x4_c, x8, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1202, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x80, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1203, x0, x1_c, x11, x12, x14_c, x15_c, x17, x19, x20_c, x21_c, x22_c, x24, x28_c, x29_c, x30_c, x31_c, x32, x34, x35, x36, x37, x39, x40_c, x41_c, x42, x44, x45, x46_c, x47_c, x48_c, x51, x52, x53_c, x56_c, x57, x58, x59_c, x62_c, x63_c, x65, x66_c, x67_c, x69_c, x70, x73, x75, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83, x84, x85_c, x87_c, x90, x91_c, x92_c, x93_c, x94, x96);
and (w1204, x6, x15, x17, x19_c, x40_c, x43, x45_c, x48, x55_c, x58_c, x62_c, x67_c, x78_c, x94);
and (w1205, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x62_c, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w1206, x73, x99_c);
and (w1207, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1208, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x77_c, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1209, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1210, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1211, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1212, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1213, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95_c, x97_c, x99_c);
and (w1214, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1215, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52, x82, x90_c, x96, x98, x99_c);
and (w1216, x4_c, x5_c, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1217, x0, x1, x3_c, x11_c, x12, x14, x19_c, x21_c, x22_c, x25_c, x27, x28, x29_c, x32_c, x33, x34_c, x35, x38, x39_c, x40, x42, x46, x47, x48_c, x50, x52_c, x54, x56, x57_c, x60, x61_c, x62_c, x63, x65_c, x66_c, x69_c, x70, x73, x76_c, x77_c, x80, x84, x88_c, x90_c, x91_c, x92_c, x93, x94_c, x97, x98);
and (w1218, x0, x1_c, x5_c, x6, x7_c, x8, x9, x10, x11, x12, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x23, x24_c, x27, x28, x29_c, x30, x32_c, x36, x37_c, x40, x41_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49, x50, x51, x52, x53_c, x54, x55, x56_c, x57_c, x58_c, x59, x62_c, x64, x65, x66, x67, x68, x69, x70, x71_c, x72_c, x73_c, x74, x77, x78, x79, x81_c, x83, x85, x86, x87_c, x88_c, x89, x90_c, x91, x93_c, x94, x95_c, x96_c, x98_c);
and (w1219, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1220, x2_c, x3, x4, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1221, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x19, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1222, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1223, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1224, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1225, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73_c, x81, x84, x85, x95, x99);
and (w1226, x0_c, x1, x2, x3, x5, x7, x9, x10_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1227, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1228, x0_c, x5, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1229, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1230, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1231, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1232, x0, x1, x2_c, x4, x5, x6, x8_c, x9, x11_c, x12_c, x13_c, x14, x17, x27_c, x29, x31, x34, x36_c, x38_c, x41, x44, x45, x48_c, x49, x50_c, x51, x52_c, x59, x63_c, x64_c, x69, x70_c, x71, x74_c, x75, x80, x83, x84_c, x85, x87, x89, x92, x97, x98, x99);
and (w1233, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92, x93_c, x97_c);
and (w1234, x0_c, x3, x4, x7_c, x8, x11_c, x12_c, x14, x30_c, x38_c, x40, x42, x49_c, x50_c, x52_c, x60_c, x73, x74, x75, x77_c, x83_c, x84, x89_c, x90, x97, x98);
and (w1235, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x32_c, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1236, x3_c, x5, x6, x7_c, x9_c, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1237, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1238, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83, x93_c, x97_c);
and (w1239, x12_c, x40, x68, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1240, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x54, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1241, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1242, x36_c, x48_c, x63_c, x80_c);
and (w1243, x6, x13_c, x21_c, x24_c, x34, x46_c, x51, x57_c, x60, x61_c, x62, x65_c, x68, x74, x92_c, x94_c);
and (w1244, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x15, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1245, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1246, x0_c, x5, x23_c, x30_c, x31, x32, x34, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1247, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1248, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x17, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1249, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1250, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89, x91_c, x92_c, x94_c);
and (w1251, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1252, x2_c, x3, x14, x15, x16, x19_c, x21_c, x22_c, x23, x24_c, x25_c, x27, x29_c, x30, x32_c, x33_c, x34, x35_c, x37, x39, x40_c, x42_c, x44_c, x47, x49_c, x55_c, x56, x60_c, x64, x66, x68_c, x69, x70, x72_c, x74_c, x76, x77_c, x78, x79_c, x82_c, x87, x88_c, x91, x92_c, x93, x95, x96, x97, x98, x99);
and (w1253, x18, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1254, x0_c, x1, x2, x3_c, x4, x5, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1255, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1256, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c);
and (w1257, x0, x2, x4_c, x6, x7_c, x9_c, x13_c, x15, x16, x19, x20, x24, x27, x29_c, x31_c, x33_c, x35, x37_c, x38_c, x39, x45_c, x50_c, x51, x52_c, x55_c, x56, x59_c, x61_c, x73_c, x76_c, x82, x89, x92_c, x95, x96_c);
and (w1258, x0, x2_c, x3, x8_c, x9, x14_c, x17_c, x18, x29_c, x32, x35, x37, x38_c, x42_c, x49, x51, x52, x57, x58_c, x59, x60_c, x68, x69, x71, x75_c, x76, x78_c, x80, x89, x90_c, x98);
and (w1259, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x20, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1260, x0_c, x5_c, x6, x12, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1261, x1_c, x2, x5_c, x7, x15_c, x17_c, x18_c, x20, x22_c, x26, x28, x36_c, x43_c, x49, x52, x55_c, x58, x59, x61, x68, x73, x75_c, x77_c, x80_c, x82, x91, x94_c, x95, x96, x98);
and (w1262, x1, x2_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1263, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1264, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x59_c, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1265, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1266, x25, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1267, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w1268, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1269, x0_c, x1_c, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1270, x1, x2_c, x6, x13_c, x14, x16_c, x17_c, x20, x21, x22, x24_c, x29_c, x31_c, x32, x34_c, x35_c, x38, x40_c, x41_c, x42_c, x47_c, x48, x49, x50_c, x52, x54, x56_c, x58_c, x60_c, x62_c, x64, x66, x70_c, x74, x76_c, x78, x79, x80_c, x83, x84, x85, x86_c, x91, x95_c);
and (w1271, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x79, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1272, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1273, x0, x1_c, x3, x4, x5_c, x7, x10, x12, x14_c, x15_c, x16, x17, x18, x20_c, x22, x23, x24_c, x25, x28, x29, x30_c, x31_c, x32, x33_c, x34_c, x35_c, x37, x38, x39_c, x40, x42_c, x43_c, x44, x46, x47, x49, x50, x51, x52_c, x57_c, x58_c, x60_c, x61, x62_c, x63_c, x65_c, x67_c, x68, x69_c, x70, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x80, x81, x82_c, x84_c, x85, x86, x87_c, x88_c, x89_c, x90, x91_c, x93_c, x94, x96, x97, x98_c);
and (w1274, x0_c, x2, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1275, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x86, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1276, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1277, x12_c, x32, x85, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1278, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49_c, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1279, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1280, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x52, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1281, x29, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1282, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x50, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1283, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x66_c, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1284, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x81_c, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1285, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1286, x5_c, x9, x27, x40, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1287, x12_c, x26_c, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1288, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1289, x13_c, x14_c, x25, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w1290, x0, x2, x3_c, x4, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16_c, x17_c, x18, x19, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x28_c, x29_c, x30, x31_c, x32, x33_c, x34_c, x35, x36_c, x37_c, x38, x39_c, x40, x41, x42, x43_c, x44, x45_c, x46, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58_c, x60, x61_c, x62_c, x63, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80, x81_c, x82, x83_c, x84_c, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91_c, x92, x93, x94_c, x96_c, x97, x98_c, x99);
and (w1291, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x50_c, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1292, x4_c, x10, x15_c, x22, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w1293, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60, x83_c);
and (w1294, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1295, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94, x95_c, x96, x98, x99);
and (w1296, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99);
and (w1297, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1298, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x61, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1299, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79, x83_c);
and (w1300, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1301, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x78_c, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1302, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1303, x5_c, x9, x27, x61_c, x76_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1304, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1305, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1306, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1307, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1308, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80_c, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1309, x8, x16, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1310, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13_c, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1311, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1312, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x52, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1313, x0_c, x2, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1314, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16_c, x83_c);
and (w1315, x0, x2, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x11_c, x12_c, x13, x14_c, x15_c, x16, x17_c, x18, x19_c, x20_c, x21, x22, x26, x27_c, x28, x29, x30, x31, x32, x34, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41, x42_c, x44, x45, x46_c, x47, x48, x49, x51_c, x52_c, x53, x55_c, x56, x58, x59, x61_c, x63, x65, x66_c, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74, x75, x76, x77_c, x78, x79_c, x80, x81, x82_c, x83, x85_c, x86, x87_c, x89_c, x92, x93, x94_c, x95_c, x96_c, x97, x98_c, x99_c);
and (w1316, x0, x1_c, x3, x4_c, x5_c, x6, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x15, x16, x17, x18, x20_c, x21_c, x22_c, x23_c, x25_c, x28, x29, x30, x31_c, x36_c, x37_c, x38_c, x39_c, x40, x41, x42, x44, x46_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55_c, x58, x61_c, x62_c, x64, x65_c, x66, x67, x69_c, x70, x72_c, x73_c, x74_c, x75_c, x76, x78_c, x79_c, x80, x81, x82, x84, x85_c, x86_c, x87_c, x88_c, x91, x92_c, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w1317, x1_c, x3, x7_c, x8, x10, x11, x13_c, x16, x17, x21_c, x24, x26_c, x35, x45_c, x48_c, x49, x50, x52_c, x53, x56, x60_c, x62_c, x63_c, x64, x66_c, x75, x78_c, x85, x86_c, x93_c);
and (w1318, x0_c, x4_c, x5, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1319, x0_c, x1_c, x2, x6, x7_c, x8, x10, x11, x12_c, x13, x14_c, x15, x17_c, x18, x19_c, x20_c, x21, x22_c, x24, x25, x26, x28, x29, x30, x31_c, x32_c, x33_c, x34_c, x36_c, x37_c, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49, x51_c, x52_c, x53_c, x54, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x69, x71_c, x72_c, x73, x75, x76_c, x77, x79_c, x80_c, x81, x83_c, x84_c, x85, x86_c, x87_c, x88_c, x89, x90, x91_c, x92, x93, x94, x95, x96_c, x97, x98_c, x99_c);
and (w1320, x0, x1, x3, x4_c, x5, x6, x7, x8_c, x9_c, x10_c, x12_c, x13_c, x14_c, x15, x16_c, x17_c, x19, x21, x22_c, x23_c, x24, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34, x35_c, x36, x38, x39_c, x41_c, x42, x43, x44_c, x45_c, x46, x47, x48_c, x51, x52, x53_c, x54_c, x55, x56, x58, x60_c, x61_c, x63, x64_c, x65, x66, x67_c, x68, x69, x70, x72_c, x73, x74_c, x75_c, x76, x77, x79, x80, x82, x83, x84_c, x85, x89_c, x90_c, x91_c, x93_c, x94_c, x95_c, x97_c, x99);
and (w1321, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x99_c);
and (w1322, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1323, x7, x14, x16, x20, x23_c, x35_c, x42_c, x43_c, x45, x58, x60_c, x64, x65, x69, x82, x85_c, x93_c, x96_c);
and (w1324, x0, x2_c, x3_c, x4_c, x5, x6, x7, x8_c, x9_c, x10_c, x11, x12_c, x15, x16, x17, x18_c, x19, x20_c, x21, x22_c, x23, x25, x26_c, x27_c, x28, x29, x30, x31, x32, x33_c, x34_c, x35, x36_c, x37, x39, x40_c, x42, x43_c, x44_c, x45, x47_c, x48_c, x49, x50_c, x52, x53_c, x54_c, x55_c, x56, x57_c, x58, x59_c, x60_c, x61, x62_c, x63_c, x64, x66, x67, x68_c, x69_c, x70_c, x71_c, x73_c, x74, x75_c, x78, x79, x80, x82, x85_c, x86_c, x87, x89_c, x90, x91_c, x93, x94, x95, x96_c, x97_c, x98, x99_c);
and (w1325, x1, x4, x11_c, x12, x14_c, x16, x17_c, x20_c, x36, x41_c, x43_c, x44_c, x46_c, x48_c, x49_c, x52, x53_c, x54, x56_c, x59, x62, x71_c, x77_c, x79_c, x80, x83_c, x86_c, x89, x90_c, x91, x95, x96);
and (w1326, x0, x1, x2, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x12_c, x13_c, x15, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28, x29, x30_c, x31, x32_c, x33_c, x34_c, x35, x36, x38_c, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50, x51, x52_c, x53_c, x55_c, x56_c, x57_c, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64, x65_c, x66_c, x67_c, x68, x70, x72_c, x73, x74_c, x78, x79, x81, x82_c, x84_c, x86, x87_c, x88, x90, x91_c, x94, x95, x97_c, x98, x99);
and (w1327, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x98_c, x99_c);
and (w1328, x12_c, x32, x52_c, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1329, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1330, x6_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1331, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x42, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1332, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x85_c, x86_c, x87, x88_c, x89, x90, x92, x94, x95, x97_c, x99_c);
and (w1333, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1334, x0, x3, x5_c, x6_c, x7_c, x9, x13, x15, x16, x20, x21_c, x24, x26_c, x27, x28, x30_c, x31, x32_c, x33_c, x35, x36, x37_c, x38, x41, x42, x43_c, x45, x46, x48_c, x49, x52, x53, x54, x56, x57_c, x58, x60_c, x61, x62_c, x64, x66, x67_c, x68_c, x70_c, x71, x72_c, x73, x75_c, x76_c, x78_c, x83, x86, x87_c, x89_c, x94, x99_c);
and (w1335, x0_c, x1, x2, x3, x4_c, x5, x6_c, x7, x9, x10_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1336, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1337, x4_c, x27, x28, x34_c, x36, x41, x53, x54_c, x57_c, x66, x68_c);
and (w1338, x1_c, x3, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x12_c, x13, x14, x15_c, x16_c, x17, x18, x20_c, x21, x22, x23, x24, x25, x26_c, x28, x30, x32_c, x33_c, x35, x36_c, x39, x40_c, x41, x44_c, x45, x47_c, x48, x49_c, x50, x54_c, x55_c, x57_c, x59, x61, x63, x64, x65_c, x66_c, x67, x69, x71, x73, x74, x75, x77_c, x79, x80, x81_c, x82, x83, x85_c, x88, x89_c, x90, x91_c, x93_c, x96, x97, x98_c, x99_c);
and (w1339, x8, x21_c, x25, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1340, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1341, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x62, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1342, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x74, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1343, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x97);
and (w1344, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x63, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1345, x5_c, x11_c, x12, x13, x15, x16_c, x18, x20_c, x21, x23, x29_c, x31_c, x37, x51, x56, x57_c, x61_c, x70, x71_c, x76, x77, x82, x89_c, x90, x92, x94);
and (w1346, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1347, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x37, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1348, x0_c, x1, x5, x6, x7, x8_c, x10, x11, x13, x18_c, x22_c, x23_c, x24, x27, x33, x34, x35_c, x40_c, x41, x42, x43, x46, x49_c, x52, x54, x56, x57_c, x59, x60, x63_c, x64_c, x66, x68, x69, x71, x72_c, x73_c, x74_c, x75_c, x77, x79, x81, x83, x84, x86_c, x87_c, x93_c, x94, x95_c, x96, x97_c, x98_c, x99_c);
and (w1349, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37_c, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1350, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x35, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1351, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1352, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x63_c, x65, x72_c, x81, x84, x85, x95, x99);
and (w1353, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x98, x99_c);
and (w1354, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x50_c, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1355, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1356, x2_c, x4, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1357, x2_c, x4, x5_c, x6, x8_c, x11_c, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1358, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15, x83_c);
and (w1359, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1360, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1361, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x32_c, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1362, x12_c, x36_c, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1363, x0, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1364, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x51, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1365, x0_c, x1, x2, x3_c, x4_c, x5, x6_c, x8_c, x9, x11_c, x12, x13, x16_c, x18, x19, x20_c, x21, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29_c, x30, x31, x32, x33, x34, x35, x36, x37_c, x38_c, x39, x40, x41, x43_c, x44_c, x45_c, x46_c, x47_c, x48, x49, x50_c, x51, x52_c, x53, x54_c, x56, x57, x58_c, x59_c, x60, x62_c, x63_c, x65, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x83, x84_c, x85_c, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92, x93, x94, x95, x96_c, x97_c, x99);
and (w1366, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c, x99_c);
and (w1367, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28, x83_c);
and (w1368, x49, x94_c, x97_c);
and (w1369, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1370, x0_c, x1_c, x4_c, x5_c, x6, x8_c, x9, x10, x12_c, x13, x14, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22_c, x23_c, x24, x26, x27, x30_c, x31_c, x33, x36, x38, x41, x42_c, x44_c, x46_c, x50_c, x51_c, x54, x55_c, x56_c, x58_c, x59_c, x60_c, x61_c, x62, x63, x64_c, x67, x68, x70, x71, x72_c, x73, x74_c, x75, x78_c, x79_c, x80, x81_c, x82, x83_c, x87, x88_c, x89, x91_c, x94, x95_c, x96_c, x97);
and (w1371, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1372, x0, x1, x2_c, x4, x6_c, x7, x8_c, x9, x10_c, x11_c, x14, x15, x16_c, x17, x18_c, x19, x20, x21_c, x22_c, x23, x24, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31_c, x32, x34_c, x35, x38, x39, x40_c, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48_c, x49, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59, x61_c, x63_c, x65_c, x67_c, x68_c, x69, x70, x72_c, x73, x75, x76, x77_c, x78_c, x79_c, x81_c, x82, x84, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99);
and (w1373, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1374, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x11_c, x12, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1375, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1376, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71, x73_c, x76, x85, x89, x93, x97_c);
and (w1377, x0_c, x2_c, x3, x4_c, x6_c, x15, x16_c, x17, x21, x23, x26, x28, x30_c, x31, x32, x35_c, x36, x37_c, x38, x39_c, x41, x43_c, x46_c, x47_c, x49, x51_c, x56_c, x59, x63_c, x64, x65, x68, x70, x75_c, x76_c, x81_c, x82, x84, x87_c, x88, x89, x90_c, x92, x99_c);
and (w1378, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x60_c, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1379, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1380, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1381, x1_c, x6_c, x14, x29_c, x49);
and (w1382, x15, x20, x21_c, x29, x41, x49_c, x58, x63_c, x64, x70, x99);
and (w1383, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x88_c, x89, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1384, x0, x1_c, x3_c, x5_c, x6, x8, x9, x10_c, x11, x12, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x23_c, x25_c, x27_c, x28_c, x29, x30_c, x31, x32_c, x34, x35, x36_c, x38, x39_c, x40_c, x41_c, x43, x44, x45, x47_c, x48_c, x50_c, x53_c, x55, x56, x58, x60, x61, x62, x64, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x74_c, x76_c, x77, x78_c, x79, x81, x82_c, x84, x85_c, x86, x87, x88, x89_c, x90, x91, x92, x93_c, x94, x95, x97_c, x98_c, x99);
and (w1385, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1386, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x55, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1387, x1_c, x9, x11, x14, x16, x22_c, x25_c, x35_c, x48_c, x55_c, x63_c, x64, x70, x75, x80_c, x85_c, x90_c, x92_c, x96_c, x97);
and (w1388, x19_c, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1389, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1390, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77_c, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1391, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1392, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1393, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1394, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35_c, x83_c);
and (w1395, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1396, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1397, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1398, x11, x12_c, x15_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1399, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1400, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1401, x0_c, x1, x2_c, x3, x4_c, x5, x6, x7_c, x8, x9, x10, x11_c, x12, x13_c, x14_c, x15, x16_c, x18_c, x19_c, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x30_c, x31_c, x32, x33, x34_c, x35, x36_c, x37_c, x38, x39_c, x40, x41_c, x42, x43, x44_c, x45, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55, x56_c, x57_c, x58, x59_c, x60_c, x61_c, x62, x63, x66, x67_c, x68, x69_c, x70, x71, x72, x74, x75_c, x76, x78, x79_c, x80, x82_c, x84, x85_c, x86_c, x87, x88, x89, x90_c, x91, x92, x93, x94, x95, x96_c, x97_c, x98_c);
and (w1402, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61_c, x73_c, x76, x85, x89, x93, x97_c);
and (w1403, x1, x2_c, x4, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1404, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1405, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x73_c, x76, x85, x89, x93, x97_c);
and (w1406, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1407, x1_c, x2, x4_c, x5, x7_c, x9, x11_c, x14_c, x15, x17, x18_c, x20_c, x21_c, x22_c, x23_c, x25, x26_c, x28, x29, x30, x31_c, x32, x33_c, x34, x36, x38, x39_c, x40, x43_c, x44_c, x47_c, x48_c, x50, x54, x58_c, x60_c, x61_c, x62, x64, x66_c, x68, x71, x73, x74, x75, x79, x81_c, x82_c, x84, x85, x88_c, x90_c, x91, x92_c, x98);
and (w1408, x16, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1409, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80_c, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1410, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71, x73_c, x76, x85, x89, x93, x97_c);
and (w1411, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1412, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1413, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43_c, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1414, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x48_c, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1415, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1416, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x74_c, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1417, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1418, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1419, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w1420, x7, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1421, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1422, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1423, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x35, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1424, x13_c, x14_c, x26, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w1425, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1426, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1427, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1428, x1, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1429, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x83, x93_c, x97_c);
and (w1430, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x87, x90, x93, x94_c, x96, x97);
and (w1431, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92_c, x94_c, x95_c, x96_c, x98, x99);
and (w1432, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1433, x2_c, x11, x29_c, x55, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1434, x2_c, x11, x29_c, x30_c, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1435, x1, x3_c, x4, x5_c, x6_c, x7_c, x9_c, x12_c, x15_c, x16, x17, x18, x19_c, x20_c, x21_c, x27, x29_c, x30_c, x32, x35_c, x39, x40, x42, x44_c, x46, x50, x51_c, x53_c, x55, x56_c, x60, x70_c, x72_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x92_c, x97_c, x99_c);
and (w1436, x4_c, x10, x15_c, x22, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1437, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93, x95, x97_c);
and (w1438, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1439, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1440, x0_c, x2, x5_c, x6, x7_c, x9_c, x10, x13_c, x14_c, x15_c, x16, x17, x18, x20, x21_c, x22_c, x23, x25_c, x26, x27, x28, x29_c, x31_c, x32_c, x33, x35_c, x36, x37_c, x38_c, x39_c, x40, x42_c, x45, x47, x48, x49_c, x51_c, x52, x55, x56, x57, x58_c, x61, x64, x67, x68, x70_c, x71, x72, x73, x74, x75, x77, x78_c, x79_c, x81, x82, x84_c, x85, x86_c, x87, x88_c, x89_c, x91_c, x92_c, x93, x94, x97);
and (w1441, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w1442, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1443, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1444, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92, x93, x94_c, x97_c);
and (w1445, x4, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1446, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36_c, x83_c);
and (w1447, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1448, x5_c, x9, x22_c, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1449, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1450, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x70, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1451, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1452, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1453, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x96, x98, x99);
and (w1454, x0, x1, x2_c, x3, x5, x6, x7, x8, x9_c, x11, x12, x13_c, x14_c, x15, x16, x17_c, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x24, x26, x28_c, x29, x30, x31, x32_c, x34, x36, x40, x41_c, x42, x46_c, x47, x49_c, x50, x52_c, x53_c, x54, x55_c, x56_c, x58, x60, x64, x65_c, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73_c, x74, x76, x78, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91_c, x92_c, x93, x94, x95_c, x96, x98, x99_c);
and (w1455, x3, x21_c, x26_c, x29, x39, x40, x55, x79, x83, x96_c, x97);
and (w1456, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1457, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1458, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87_c, x93_c, x97_c);
and (w1459, x0, x3, x10, x12, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1460, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x90_c, x91, x93, x95_c, x96, x98, x99);
and (w1461, x13_c, x14_c, x37_c, x39_c, x44, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1462, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1463, x27, x28_c, x29_c, x34, x45_c, x46, x48, x52_c, x62_c, x82_c, x95, x99_c);
and (w1464, x0_c, x3, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w1465, x17, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1466, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86, x89, x93, x97_c);
and (w1467, x6_c, x7, x8_c, x12_c, x13_c, x14, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1468, x21_c, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1469, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1470, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x32_c, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w1471, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1472, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1473, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1474, x1_c, x2, x3, x4, x5_c, x6_c, x8, x12_c, x13, x14_c, x15, x16, x17, x18, x20, x21, x23, x27, x29, x30_c, x31, x34, x36, x37, x41_c, x42_c, x44_c, x45, x46_c, x48, x49, x50_c, x51_c, x53_c, x55, x56, x59_c, x61_c, x62_c, x63, x64, x65, x66_c, x69_c, x73_c, x74_c, x75, x76, x77, x80_c, x82_c, x83, x85_c, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x94_c, x97, x98);
and (w1475, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1476, x0, x3, x10, x13, x14, x15, x16_c, x22, x28, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1477, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1478, x6, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1479, x3_c, x5_c, x6, x7_c, x8_c, x10, x11_c, x12, x13_c, x14_c, x15, x16_c, x17, x18_c, x19_c, x22_c, x23, x24, x25_c, x27_c, x28, x29_c, x31, x33, x34, x35, x36_c, x38_c, x39, x40, x41_c, x42_c, x43_c, x44, x45_c, x46, x47_c, x49, x50_c, x51, x53, x54_c, x55, x57, x58_c, x59_c, x61_c, x62, x63, x64_c, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x71, x72, x74, x75_c, x76, x78, x79, x80, x81_c, x82_c, x84, x85, x86_c, x87, x88, x89_c, x90_c, x92_c, x93_c, x96, x98, x99);
and (w1480, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w1481, x0_c, x1, x2, x3_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
assign w1482 = x23_c;
and (w1483, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1484, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1485, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x91_c, x93_c, x94_c, x96_c, x97, x98, x99_c);
and (w1486, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1487, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x77_c, x82, x83, x93_c, x97_c);
and (w1488, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1489, x0, x1, x2_c, x3, x4_c, x5_c, x6_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1490, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1491, x12_c, x32, x80, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1492, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x35_c, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1493, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x63, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1494, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x58_c, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1495, x3_c, x5, x7_c, x8, x9, x10, x11, x13_c, x18, x20, x21_c, x22, x23_c, x24, x27_c, x28, x29_c, x31, x33_c, x36, x37_c, x41, x42_c, x46, x49_c, x50, x51, x56_c, x58, x59, x60, x61, x64, x67, x68, x69, x71, x72, x74_c, x75, x77, x78_c, x79, x81, x86_c, x87_c, x89_c, x91, x95, x96_c, x97);
and (w1496, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1497, x0, x1_c, x2_c, x3_c, x4_c, x5, x6, x7_c, x8_c, x9_c, x10, x11_c, x12_c, x13, x14_c, x15, x16, x17_c, x18_c, x19_c, x20, x21, x22_c, x23, x24_c, x25_c, x26, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x34, x35_c, x36, x37_c, x38_c, x40, x41_c, x42, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51_c, x52, x53, x54_c, x55_c, x56_c, x57_c, x58_c, x59, x60, x61, x62, x63, x64, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75, x76_c, x77, x78, x79, x81, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1498, x3_c, x18, x27_c, x34_c, x73_c, x98);
and (w1499, x0, x1, x2, x3_c, x4, x5_c, x6, x7_c, x8_c, x9_c, x10, x11_c, x12, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27, x28_c, x29_c, x30, x31_c, x32, x33_c, x34, x35, x36_c, x37_c, x38, x39, x40_c, x41, x42_c, x43, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50_c, x51, x52_c, x53_c, x54, x55, x56, x57, x58_c, x59, x60, x61, x62, x63, x64, x65, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x73, x74_c, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97_c, x98, x99);
and (w1500, x12_c, x40, x44_c, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1501, x0_c, x2_c, x5, x7, x8_c, x11, x13, x14_c, x16, x18_c, x19, x20, x21_c, x22, x23, x24_c, x25, x26_c, x27, x29_c, x35_c, x36_c, x40_c, x42, x46_c, x48_c, x49, x58, x59, x60, x61, x62, x63, x64, x65_c, x66_c, x67, x68_c, x69_c, x70_c, x75_c, x76_c, x77_c, x79_c, x82_c, x83, x84_c, x87, x88, x90_c, x91, x92, x93, x94_c, x98);
and (w1502, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x83, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1503, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x95, x98_c, x99_c);
and (w1504, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x70_c, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1505, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1506, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1507, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92, x95, x97, x98, x99_c);
and (w1508, x0, x1_c, x2, x3_c, x4, x5_c, x6, x7_c, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27_c, x28, x29, x31_c, x32_c, x34_c, x35_c, x36, x38, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x47_c, x48, x49_c, x51, x52_c, x54_c, x55, x57, x58_c, x59_c, x60, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69, x70, x71_c, x73, x74, x75, x76, x77_c, x78, x79_c, x80, x81_c, x82_c, x83, x84_c, x85_c, x87_c, x88_c, x90_c, x91, x93, x95, x96, x97, x98_c, x99);
and (w1509, x6, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1510, x0, x5_c, x7, x13, x14_c, x15, x16_c, x19_c, x23, x24, x25_c, x27, x28, x29, x36, x37_c, x39_c, x40_c, x41, x43, x50_c, x51, x55_c, x57_c, x63_c, x64_c, x67_c, x69_c, x73_c, x74, x76_c, x82_c, x90, x91_c, x95, x96);
and (w1511, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x37, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1512, x0, x2_c, x5_c, x9, x10, x13, x15, x18, x22, x26_c, x29, x30, x31, x33, x35_c, x39, x40_c, x41, x42, x45, x46, x48_c, x49_c, x52_c, x57_c, x59, x60, x62_c, x63_c, x66, x69, x70_c, x72, x73, x74_c, x75, x79, x81, x87, x90, x91, x92, x93, x94_c, x96_c);
and (w1513, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1514, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1515, x2_c, x11, x29_c, x96_c, x98, x99);
and (w1516, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1517, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1518, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x68_c, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1519, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1520, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x42, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1521, x1, x2, x3, x5_c, x6_c, x9, x12_c, x13, x14_c, x15, x16, x17_c, x18_c, x19, x20, x21, x24, x26, x27, x28, x29, x30_c, x31, x34_c, x35_c, x36_c, x37_c, x43, x45_c, x46, x47, x49, x50_c, x51, x52, x53_c, x56, x58, x61_c, x62, x65_c, x69_c, x70, x71, x72, x74_c, x75, x76, x77, x78, x81_c, x82, x83_c, x88, x90, x91_c, x92_c, x96_c, x97_c, x98, x99_c);
and (w1522, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1523, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91, x92, x93_c, x95, x96_c, x98, x99_c);
and (w1524, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1525, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1526, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1527, x12_c, x32, x77, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1528, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1529, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x17, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1530, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1531, x0, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1532, x4_c, x10, x15_c, x22_c, x24, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1533, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1534, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1535, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x30, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1536, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1537, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x88_c, x89, x90_c, x92_c, x93, x95_c);
and (w1538, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x88_c, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1539, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x50, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1540, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1541, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1542, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1543, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1544, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1545, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1546, x1_c, x2, x3, x4, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x13_c, x14, x15_c, x16, x17_c, x18_c, x19_c, x20, x21_c, x22_c, x23, x24_c, x25_c, x27_c, x28, x29, x30, x31_c, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50_c, x51_c, x52_c, x54, x55_c, x56_c, x57_c, x58_c, x59, x60_c, x61, x62, x64, x66_c, x67, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76, x77, x78_c, x79, x81_c, x82_c, x83_c, x84, x85, x86_c, x87, x88, x89, x90_c, x91, x92_c, x93_c, x94_c, x95, x96, x97, x98_c, x99_c);
and (w1547, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1548, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1549, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1550, x33, x34_c, x36_c, x40, x41_c, x63, x66_c, x67, x71_c, x94_c, x97_c);
and (w1551, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1552, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1553, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x36, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1554, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1555, x0, x1, x2, x3_c, x4_c, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20_c, x21_c, x22, x23_c, x25, x26, x27, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35, x36_c, x37, x39, x40_c, x41_c, x42, x43, x44_c, x46_c, x47, x48, x49, x50, x51, x52_c, x53_c, x54, x55, x56_c, x57_c, x58_c, x59, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70, x71_c, x74_c, x76_c, x77_c, x78, x79_c, x80_c, x81, x82, x83, x84_c, x86, x87_c, x88_c, x89_c, x90, x91_c, x92, x93, x94, x95, x98, x99_c);
and (w1556, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x65_c, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1557, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1558, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95, x96, x98, x99_c);
and (w1559, x0_c, x2_c, x5_c, x7_c, x8_c, x9, x10, x11_c, x13_c, x14_c, x20, x21_c, x23, x24, x25_c, x26, x27, x28_c, x29_c, x30, x32, x33, x36, x37, x38, x39, x40, x45_c, x49, x50, x53_c, x54_c, x55_c, x57, x58_c, x60_c, x61, x62_c, x63_c, x64, x72_c, x73_c, x77_c, x78_c, x80_c, x81_c, x84, x86, x87_c, x91, x92, x93_c, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w1560, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x79_c, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1561, x0_c, x4_c, x5_c, x6_c, x8, x13_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1562, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1563, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98);
and (w1564, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x97_c);
and (w1565, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x77, x79, x90_c, x93_c, x97_c);
and (w1566, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x48_c, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1567, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91, x92, x93_c, x94_c, x95, x96_c, x98, x99);
and (w1568, x0_c, x2, x3, x4, x5, x6, x7, x10_c, x11, x12, x13, x14_c, x15_c, x16_c, x17_c, x18, x19_c, x21, x23_c, x24, x25_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36_c, x37, x38_c, x39, x40, x42, x43_c, x44, x45, x46, x48_c, x49, x50, x51, x52, x53, x54, x55_c, x57, x58_c, x59_c, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70, x71, x72, x74_c, x76_c, x77, x78, x79, x80_c, x81_c, x83, x84, x85_c, x86, x88, x89_c, x90, x91, x92, x93, x94, x95_c, x96, x97_c, x98, x99);
and (w1569, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1570, x5, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1571, x0_c, x1, x2, x3, x4_c, x5_c, x6, x7_c, x8_c, x9_c, x11, x12, x14_c, x15, x16_c, x17, x18, x20_c, x21_c, x22, x23, x25_c, x27_c, x28, x29_c, x30_c, x31, x32, x33_c, x34_c, x35_c, x36_c, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46, x47, x48, x49_c, x50, x51, x52_c, x53_c, x54_c, x55, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64_c, x67_c, x68, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76, x79, x81_c, x82_c, x83_c, x84_c, x85, x86, x87_c, x88_c, x89, x90, x91_c, x93_c, x94, x95_c, x96_c, x97, x98_c);
and (w1572, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x58_c, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1573, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1574, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1575, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1576, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x95, x96, x97_c);
and (w1577, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84, x93_c, x97_c);
and (w1578, x12_c, x32, x78, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1579, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x71, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1580, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1581, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1582, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x76_c, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1583, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x98_c, x99_c);
and (w1584, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1585, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x60, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1586, x1, x2_c, x6, x7_c, x8, x9, x10, x11, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1587, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1588, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x12, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1589, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x76, x85, x89, x93, x97_c);
and (w1590, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1591, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x29_c, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1592, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x82, x90_c, x96, x98, x99_c);
and (w1593, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x7, x9_c, x10_c, x14, x16_c, x18, x19_c, x20, x21, x23, x24, x25_c, x26_c, x27, x28_c, x29, x30, x31_c, x32, x33_c, x34_c, x35, x36, x37_c, x38_c, x40, x41_c, x44_c, x45, x46_c, x50_c, x51, x52_c, x53_c, x54, x55_c, x56_c, x57, x58, x59, x61, x62, x63, x64_c, x66, x67, x68, x69, x71_c, x72_c, x73, x75_c, x77, x79, x80_c, x81, x82, x83, x84, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93, x98_c);
and (w1594, x3_c, x5, x7, x8_c, x14, x15_c, x17_c, x21_c, x27_c, x31, x35, x38_c, x39_c, x41, x44_c, x45_c, x47_c, x51_c, x55_c, x58_c, x59_c, x64_c, x66_c, x67_c, x69_c, x76_c, x81_c, x82_c, x85, x99);
and (w1595, x0, x1, x2_c, x3, x4, x6, x7_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1596, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x96, x97, x98, x99_c);
and (w1597, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1598, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1599, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x94, x95, x97_c, x99_c);
and (w1600, x8, x9_c, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1601, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1602, x0, x1, x2_c, x5_c, x7, x8_c, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18_c, x19_c, x20, x21_c, x22, x23, x24, x26_c, x27_c, x29_c, x30_c, x31, x32_c, x34_c, x35_c, x36, x37_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x46, x47, x48_c, x49, x51_c, x52_c, x53, x54, x55_c, x56_c, x57, x58_c, x59_c, x60_c, x61_c, x62_c, x63_c, x64, x65, x66_c, x67, x68_c, x69, x70_c, x71_c, x72, x73, x74, x75, x76, x77, x78_c, x79_c, x82_c, x83, x84, x85, x86_c, x87, x88, x89, x90, x91, x94_c, x95_c, x96, x97_c);
and (w1603, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91, x93_c, x95_c, x96, x98, x99);
and (w1604, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1605, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1606, x9, x10_c, x16_c, x20_c, x44, x47, x52, x60_c, x76, x84_c);
and (w1607, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1608, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1609, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54, x83_c);
and (w1610, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1611, x12_c, x40, x73_c, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1612, x12_c, x34, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1613, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1614, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1615, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21, x83_c);
and (w1616, x0, x1_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1617, x0_c, x4_c, x5_c, x6_c, x8_c, x9_c, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1618, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x77_c, x79_c, x82, x90, x93_c, x97_c);
and (w1619, x0_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1620, x12_c, x24, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1621, x1, x14_c, x26_c);
and (w1622, x0, x5, x6_c, x7, x9_c, x10_c, x12_c, x14, x15_c, x16_c, x17_c, x18, x20, x21, x22, x25, x26_c, x27_c, x29, x30_c, x32_c, x33, x34_c, x36, x37_c, x38, x39, x40, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x52_c, x53, x54, x55_c, x56_c, x57, x59, x60_c, x61_c, x63_c, x64_c, x65_c, x66, x67, x68, x69_c, x70, x71_c, x74_c, x75_c, x76, x77, x78, x79, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86, x87_c, x88, x89, x91, x92, x95_c, x96_c, x98_c, x99);
and (w1623, x0_c, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1624, x0_c, x4_c, x5, x12_c, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1625, x11, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1626, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1627, x8_c, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1628, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x95, x96_c, x98, x99_c);
and (w1629, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x38, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1630, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x72, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1631, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1632, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1633, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1634, x0_c, x1, x3_c, x5_c, x6, x7, x9_c, x10_c, x11, x12_c, x14, x16_c, x17_c, x22_c, x23, x26_c, x28_c, x29, x32_c, x33, x35_c, x36_c, x38, x39_c, x40_c, x41_c, x43, x44, x46_c, x49_c, x50, x54, x55_c, x57, x64_c, x67_c, x71_c, x73, x74, x75_c, x76, x78, x79, x81_c, x82, x84, x86, x87_c, x89_c, x91, x93_c, x96, x99_c);
and (w1635, x12_c, x40, x55, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1636, x0_c, x5, x17, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1637, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43_c, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1638, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x84, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1639, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1640, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x85_c, x86_c, x87, x88_c, x89, x90, x92, x95, x96, x97_c, x98_c, x99_c);
and (w1641, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x62, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1642, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1643, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1644, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1645, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x19, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1646, x0, x1, x2, x5_c, x9, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1647, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x85_c, x89, x93, x97_c);
and (w1648, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x53, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1649, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91, x92, x93_c, x94_c, x95, x96, x97, x98_c);
and (w1650, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x42, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1651, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x98, x99_c);
and (w1652, x0_c, x5_c, x6, x10_c, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1653, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1654, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1655, x0_c, x1, x3_c, x5, x6_c, x8, x9, x10, x17_c, x18, x20_c, x21_c, x22, x24_c, x30, x31, x32, x33, x34_c, x37_c, x38_c, x42, x46, x47_c, x50, x53_c, x54_c, x55, x58, x59, x60, x61, x62, x63, x65, x66_c, x67, x69, x70, x71_c, x72, x73_c, x74, x75_c, x85, x87, x90, x91_c, x98_c, x99_c);
and (w1656, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x83_c, x93_c, x97_c);
and (w1657, x2_c, x4_c, x10, x16, x20, x21, x22_c, x29, x31_c, x32, x40, x45, x47, x50, x53_c, x55, x56, x57_c, x59_c, x61_c, x63, x65_c, x66_c, x70_c, x73, x74, x75, x78_c, x80_c, x87_c, x88, x98, x99);
and (w1658, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1659, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x36, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1660, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1661, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1662, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1663, x0, x1, x2, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14_c, x15_c, x16, x17_c, x18, x19_c, x20, x21, x22, x23, x24, x25_c, x26_c, x27, x28, x29_c, x30, x31, x32, x33_c, x34, x35, x36, x37_c, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46, x47, x48_c, x49, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x67, x68_c, x69_c, x70, x71_c, x73_c, x74_c, x75, x76_c, x77, x78_c, x79_c, x80_c, x81, x82, x83_c, x84, x85, x86_c, x87_c, x88_c, x89, x90, x91_c, x92, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w1664, x0, x2, x5, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1665, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1666, x0, x2, x11_c, x19_c, x20_c, x30_c, x34_c, x37_c, x40_c, x54, x57_c, x62_c, x78, x79, x80_c, x95, x99_c);
and (w1667, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1668, x11, x12_c, x15, x17_c, x21_c, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1669, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1670, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1671, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1672, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1673, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1674, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w1675, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1676, x0, x1_c, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1677, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1678, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1679, x3, x9, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1680, x0, x3, x10, x13, x14, x15, x16_c, x22, x25, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1681, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97, x99);
and (w1682, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1683, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1684, x49, x72, x73_c, x74_c, x79, x90_c, x93_c, x97_c);
and (w1685, x5, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1686, x12_c, x40, x53_c, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1687, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1688, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x13_c, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1689, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1690, x20_c, x25_c, x32, x53, x55_c, x57_c, x77_c, x79_c);
and (w1691, x4_c, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1692, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1693, x8, x21_c, x25_c, x27_c, x34, x36, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1694, x12_c, x26, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1695, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1696, x1, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1697, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1698, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x80, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1699, x0, x2, x5, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1700, x22_c, x24_c, x33_c, x37, x43_c, x53, x63, x65, x76, x90_c, x92_c, x96, x99);
and (w1701, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x49_c, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1702, x0_c, x2_c, x6_c, x7_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w1703, x6_c, x9_c, x11, x15, x16_c, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w1704, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x50, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1705, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1706, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1707, x0, x1_c, x2_c, x4_c, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w1708, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1709, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1710, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1711, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x49, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1712, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1713, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1714, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x92_c, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1715, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x52, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1716, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1717, x49, x54, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1718, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x27, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1719, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47_c, x83_c);
and (w1720, x0, x1, x2, x3, x4, x5_c, x6_c, x7, x8, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x23_c, x24, x25_c, x26, x27, x30, x31, x32_c, x33, x34, x36, x38, x39_c, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48_c, x49_c, x50, x51_c, x52, x53, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62, x63_c, x64_c, x65, x67_c, x68, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78, x80, x81, x82, x83_c, x84, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95_c, x96_c, x97_c, x98, x99);
and (w1721, x13_c, x49, x64, x69_c, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w1722, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1723, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90, x91_c, x92_c, x93_c, x96, x97_c);
and (w1724, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x25_c, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1725, x5, x10, x16_c, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1726, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x89, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1727, x1, x2_c, x3, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1728, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x38_c, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1729, x0, x2_c, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1730, x3, x5_c, x6_c, x7_c, x9, x11_c, x12, x14_c, x15_c, x18, x19_c, x20, x21, x22_c, x25_c, x29_c, x30_c, x38, x39_c, x41, x44_c, x46, x47, x48_c, x50_c, x52_c, x53_c, x55_c, x57, x58, x59, x61_c, x62_c, x63_c, x70, x73_c, x74_c, x78_c, x82, x85_c, x86_c, x87_c, x88, x90, x92, x95, x96_c, x97, x98_c);
and (w1731, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46_c, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1732, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x54_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1733, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46, x83_c);
and (w1734, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x90, x91, x92, x95, x97_c);
assign w1735 = x89_c;
and (w1736, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1737, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1738, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x86_c, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1739, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82_c, x90_c, x93_c, x97_c);
and (w1740, x5_c, x9, x27, x61_c, x69, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1741, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x71_c, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1742, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x63, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1743, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x12_c, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1744, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1745, x0, x1_c, x2_c, x3, x4_c, x5, x7, x8_c, x10, x12, x13_c, x14, x16_c, x17, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x43, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x55, x56_c, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x67, x68_c, x70_c, x71, x72, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x80_c, x81_c, x82, x83, x84, x85, x86_c, x88, x89, x90_c, x91, x92_c, x93, x94_c, x95, x96_c, x97, x98, x99);
and (w1746, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1747, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w1748, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1749, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x39_c, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1750, x49, x67_c, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1751, x0, x1, x2, x3, x5, x6, x7, x8, x9_c, x10_c, x11, x13_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19, x20_c, x23_c, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31, x33_c, x34_c, x35_c, x36_c, x37, x38, x39_c, x40_c, x42, x43_c, x44, x45, x46_c, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x57, x58_c, x59_c, x60_c, x61_c, x62_c, x64_c, x65_c, x67_c, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77, x78, x79_c, x80_c, x81, x82_c, x84, x85_c, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94, x95, x96_c, x98, x99_c);
and (w1752, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1753, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x41, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1754, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61_c, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1755, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x46, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1756, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1757, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x77_c, x79_c, x82_c, x90_c, x93_c, x97_c);
and (w1758, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x92_c, x93_c, x94, x95, x96, x97);
and (w1759, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x75_c, x77, x81_c, x82_c, x88_c, x93_c, x95_c);
and (w1760, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35_c, x40, x82, x90_c, x96, x98, x99_c);
and (w1761, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1762, x1, x3, x4_c, x8_c, x9, x10_c, x13, x15_c, x16_c, x18_c, x19_c, x20_c, x23_c, x24_c, x25_c, x26_c, x27_c, x29_c, x31, x33_c, x36_c, x37_c, x38_c, x40, x43_c, x45_c, x46, x47, x48, x49_c, x51, x52_c, x53, x54_c, x55_c, x56, x61, x62_c, x63_c, x65, x66_c, x67, x68_c, x71_c, x72_c, x73_c, x75, x76_c, x77_c, x78, x79_c, x80_c, x82, x83, x84, x85, x86_c, x87, x88, x90_c, x91, x92_c, x93, x94, x95, x96, x97, x98);
and (w1763, x0_c, x1, x2, x6, x7_c, x8_c, x9, x10, x11_c, x12, x14_c, x15, x16_c, x18, x20, x22_c, x23_c, x24_c, x25_c, x26, x27, x31_c, x33, x34, x35, x36, x38_c, x40_c, x41_c, x42, x43_c, x44, x45_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x55, x57_c, x58, x59, x60_c, x61_c, x62, x64, x65, x66, x67, x68_c, x70_c, x73, x74, x75, x76_c, x77, x78, x80, x81, x82_c, x83_c, x84_c, x86_c, x87_c, x89, x90_c, x91_c, x92_c, x94, x95_c, x96, x97_c, x99_c);
and (w1764, x0_c, x5, x23_c, x30_c, x31_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1765, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1766, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1767, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x72, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1768, x5, x12_c, x16, x31, x44, x52, x53, x61, x73_c, x74, x75_c, x77, x78_c, x81, x82_c, x84, x87, x90);
and (w1769, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31, x40, x82, x90_c, x96, x98, x99_c);
and (w1770, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x77, x82, x83, x93_c, x97_c);
and (w1771, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1772, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x61, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1773, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1774, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1775, x0, x3, x10, x13, x14, x15, x16_c, x21_c, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1776, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1777, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1778, x0, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x11, x12, x13_c, x15_c, x17, x18, x20_c, x21_c, x22_c, x23_c, x24_c, x25, x28_c, x29_c, x31_c, x32, x33_c, x34_c, x35, x36_c, x37, x38, x39, x40_c, x42, x43_c, x44, x45_c, x46_c, x47, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x58_c, x59, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70, x72, x73_c, x75_c, x76, x80, x81_c, x82_c, x84_c, x85, x88_c, x89_c, x91_c, x94_c, x95, x96, x97);
and (w1779, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x85, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1780, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1781, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50_c, x83_c);
and (w1782, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1783, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1784, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1785, x0, x2, x4, x15_c, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1786, x0, x1_c, x2_c, x3_c, x4, x5, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23_c, x25, x26, x27, x28_c, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39, x40, x42, x43, x44_c, x45_c, x46_c, x47, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x65_c, x66_c, x67, x68_c, x70, x71, x72_c, x73, x74, x75, x76_c, x77_c, x79_c, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88, x89_c, x90, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1787, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1788, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x15, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1789, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x36, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1790, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x90_c, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1791, x0_c, x1, x3, x4, x5, x7, x9, x10_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1792, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30_c, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1793, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1794, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1795, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x84, x90_c, x96, x98, x99_c);
and (w1796, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x17, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1797, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87, x93_c, x97_c);
and (w1798, x0_c, x1_c, x2, x3_c, x4, x6, x7_c, x8, x9, x10_c, x12_c, x13_c, x14, x15, x16, x17_c, x18, x19, x20, x21, x23, x24_c, x25_c, x26_c, x28_c, x29_c, x30, x32, x33, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x47_c, x48_c, x50, x51, x52, x53, x54, x55, x56_c, x57_c, x58, x59_c, x60, x61_c, x62_c, x63, x64_c, x65, x66, x68, x69, x70, x71, x72_c, x73, x74_c, x75_c, x76_c, x77, x78_c, x79, x80, x81, x82, x83, x84_c, x86, x87_c, x88_c, x89, x90_c, x91, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w1799, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1800, x1, x5, x12_c, x19_c, x30, x38_c, x45_c, x47, x48, x49_c, x50, x52_c, x54, x57_c, x60, x73_c, x77, x80_c, x82_c, x88, x96, x97);
and (w1801, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1802, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x11_c, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1803, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x71, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1804, x0_c, x1_c, x2, x3_c, x4, x5_c, x6_c, x7_c, x8, x9, x10, x11_c, x12_c, x13, x14_c, x15, x16_c, x17_c, x18, x19_c, x20, x21_c, x22_c, x23_c, x24_c, x25, x27_c, x28, x29, x30_c, x31, x32_c, x33, x34, x36_c, x37, x38, x39_c, x40, x41_c, x42, x43, x44, x45, x46_c, x47_c, x48_c, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56, x57_c, x58_c, x59_c, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x67, x68_c, x69, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80, x81_c, x82_c, x83, x84, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91, x92_c, x93, x94, x95, x96, x97, x98_c, x99_c);
and (w1805, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1806, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1807, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x38, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1808, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x28_c, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1809, x0_c, x2_c, x6_c, x7, x8, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w1810, x0_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1811, x2_c, x3_c, x4, x6, x9, x11_c, x12, x13, x14_c, x15, x16_c, x18, x19_c, x20_c, x22_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x31, x32, x34, x35, x36_c, x37, x38_c, x39_c, x41_c, x43, x45, x46_c, x49, x50_c, x51_c, x52_c, x54, x55, x56_c, x58, x60_c, x62_c, x63_c, x64, x66_c, x67_c, x69_c, x70, x71_c, x74, x76_c, x77_c, x78, x81, x82_c, x83, x84_c, x85_c, x86, x87_c, x89, x90, x91, x92, x93, x94_c, x95_c, x96, x97_c, x99);
and (w1812, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x87, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w1813, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x78, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1814, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w1815, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1816, x0, x1, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1817, x0_c, x2, x3, x4_c, x5, x8_c, x10, x11, x12, x13, x14_c, x15_c, x17_c, x18, x19_c, x20, x21, x22, x23, x24_c, x25_c, x27_c, x29, x30_c, x31, x33, x34, x35, x36, x37, x38, x40_c, x41_c, x42, x43, x44_c, x45, x46_c, x47_c, x49_c, x50, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x61_c, x62, x63, x65_c, x66, x67, x68, x69, x70, x72, x73, x74_c, x75, x76_c, x78_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x87_c, x88_c, x90, x91, x92_c, x93, x94, x95_c, x97);
and (w1818, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1819, x1_c, x2, x4, x5, x11, x12_c, x15, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1820, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1821, x9_c, x17_c, x26, x27, x28, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1822, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x29, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1823, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1824, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97, x98, x99_c);
and (w1825, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x95, x96, x97, x99_c);
and (w1826, x0_c, x1_c, x2, x4, x6, x10, x11, x12_c, x13, x14, x15, x16, x17, x19, x20, x21_c, x22_c, x23, x24, x26_c, x27_c, x30_c, x31_c, x32, x34_c, x35, x37_c, x43_c, x47_c, x48_c, x49, x50_c, x51_c, x52_c, x53, x54, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x64, x65, x66, x69_c, x71, x72, x75, x77_c, x79, x81_c, x82, x83_c, x84_c, x85, x86, x88_c, x90, x91_c, x92_c, x93_c, x95_c, x96_c, x97, x98_c, x99);
and (w1827, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1828, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1829, x2_c, x6, x8_c, x12_c, x13_c, x15_c, x16_c, x18_c, x24, x26_c, x31_c, x34, x35_c, x52_c, x56_c, x62, x64, x69, x75, x77, x88_c, x89_c, x95);
and (w1830, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x76_c, x85, x89, x93, x97_c);
and (w1831, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x45_c, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1832, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x34_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1833, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x91_c, x92, x95, x97_c);
and (w1834, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x89, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1835, x8, x21_c, x25_c, x27_c, x34, x37_c, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1836, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44_c, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1837, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x71, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1838, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1839, x4_c, x5_c, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1840, x0, x1, x2, x3_c, x4_c, x5, x6, x9_c, x10_c, x12_c, x13_c, x14_c, x15_c, x17, x19, x20, x21, x22, x23_c, x24_c, x26, x27_c, x29, x30, x31_c, x33, x34, x36_c, x37_c, x40_c, x43_c, x45_c, x46_c, x47_c, x49, x50_c, x54_c, x55_c, x56, x57, x59_c, x60_c, x61_c, x62, x64, x65, x67, x69_c, x70, x73_c, x74_c, x75_c, x78, x79_c, x80, x81_c, x82_c, x83, x84, x86_c, x87, x88_c, x89_c, x92, x93, x95_c, x96_c, x97);
and (w1841, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92_c, x95, x96, x97, x99_c);
and (w1842, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1843, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x90_c, x93, x95, x96, x97, x99_c);
and (w1844, x0, x2, x3, x6_c, x10_c, x11, x13_c, x20, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1845, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48_c, x82, x90_c, x96, x98, x99_c);
and (w1846, x0, x1_c, x3_c, x4, x7, x8_c, x10, x12_c, x13, x15, x17, x18, x19_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27, x29, x30_c, x32_c, x34_c, x37_c, x38, x40_c, x41, x42_c, x43, x47_c, x50_c, x51, x52, x53, x54, x55_c, x57_c, x58, x59_c, x61, x62, x63, x65, x66, x67, x69_c, x70_c, x71, x72_c, x73, x74_c, x75, x76, x78_c, x79, x81_c, x83, x86_c, x88_c, x89_c, x90_c, x91_c, x97, x98_c);
and (w1847, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1848, x1, x2_c, x3_c, x4_c, x5_c, x6, x8_c, x11_c, x12, x13, x14_c, x15, x17_c, x20, x21, x22, x24_c, x26, x28, x29_c, x30_c, x31, x32, x33, x34_c, x35, x36_c, x38, x39_c, x40, x41_c, x42, x43_c, x44, x45, x47, x48, x49_c, x50, x51_c, x53_c, x54, x55, x56, x57, x58_c, x60_c, x61_c, x62_c, x63, x64_c, x66_c, x67, x68, x72_c, x73, x74, x75_c, x76_c, x77, x78, x79_c, x80, x82, x84, x85, x86_c, x87_c, x91_c, x92, x93_c, x94_c, x96, x97_c, x98, x99);
and (w1849, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x46_c, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1850, x1, x2_c, x3_c, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1851, x0_c, x2, x3, x5_c, x6_c, x7, x9, x10, x11_c, x12_c, x13_c, x14_c, x17, x18_c, x20_c, x23_c, x25, x26, x27_c, x29, x30, x31_c, x36_c, x37, x38_c, x39, x40, x41_c, x42, x43_c, x44_c, x46, x47, x48, x49, x50_c, x51, x52_c, x53_c, x54_c, x56, x57_c, x58_c, x60, x61, x62, x63_c, x64, x65_c, x66, x67, x70_c, x72, x74, x75_c, x77, x78_c, x79_c, x81, x82_c, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90, x91_c, x92, x96, x97_c, x99);
and (w1852, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x87_c, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1853, x11_c, x15_c, x16, x18, x21, x23, x71_c);
and (w1854, x41_c, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1855, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x49, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1856, x0_c, x1_c, x2, x3, x8, x9_c, x12_c, x13_c, x14_c, x15_c, x18_c, x19, x20_c, x24_c, x26_c, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35, x37_c, x38_c, x39, x41, x44, x45_c, x46_c, x48, x49_c, x52, x53, x60_c, x62_c, x63, x67_c, x70, x71, x74_c, x75, x76, x78_c, x80_c, x83_c, x84, x86, x88_c, x93_c, x95);
and (w1857, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x58, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1858, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x78, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1859, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1860, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1861, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x9_c, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1862, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1863, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x49, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1864, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1865, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1866, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1867, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1868, x2_c, x4_c, x8_c, x9, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1869, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1870, x0_c, x1_c, x2_c, x3, x4, x5_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1871, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x77, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1872, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x23, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1873, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1874, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x86, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1875, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1876, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x31, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1877, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x62_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1878, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c, x99);
and (w1879, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1880, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x45, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1881, x13_c, x14_c, x22_c, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w1882, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x38_c, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1883, x8, x32_c, x57, x76_c, x79_c, x97_c);
and (w1884, x0, x2_c, x3_c, x4, x6_c, x7, x8, x11, x12, x13, x14, x17, x19_c, x20_c, x21_c, x22_c, x23_c, x24, x25, x27, x28_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x37_c, x38_c, x41_c, x42_c, x43, x44, x46, x47_c, x50, x54, x55_c, x56_c, x57_c, x58_c, x59_c, x61, x62_c, x63_c, x64_c, x66, x67_c, x68, x69_c, x70_c, x71_c, x72, x73_c, x74_c, x75_c, x77_c, x78, x79_c, x80, x82, x83, x84_c, x85_c, x86, x87_c, x88, x90_c, x91_c, x95, x96, x98_c, x99);
and (w1885, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x74, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1886, x0_c, x5, x23_c, x30_c, x31, x32, x37, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1887, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1888, x13_c, x14_c, x37, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1889, x0, x1, x3_c, x4, x5, x7, x10_c, x13, x14, x15, x17, x18_c, x19, x22, x23_c, x24_c, x28_c, x30, x32_c, x33_c, x37_c, x38, x40, x41, x44_c, x46, x47_c, x53, x57_c, x59_c, x68_c, x71, x74_c, x75, x77_c, x78, x79, x82, x83_c, x89, x90_c, x93, x96_c, x97_c);
and (w1890, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x25, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1891, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1892, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w1893, x0, x4, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x12, x13, x14, x16_c, x17, x19_c, x20, x21_c, x22_c, x23, x24, x26_c, x27, x29_c, x30, x31_c, x33_c, x34_c, x35, x36_c, x37_c, x38, x39_c, x40, x41, x43_c, x44, x46, x48, x49, x50, x51, x52, x53_c, x54_c, x55, x56, x57, x58, x60_c, x63, x64_c, x65, x66_c, x67_c, x68, x70, x71, x72, x73, x74, x75_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84, x88, x89_c, x90_c, x91_c, x92, x94, x95_c, x96_c, x97, x99_c);
and (w1894, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1895, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79, x83_c);
and (w1896, x0_c, x1, x2, x3_c, x4, x5_c, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1897, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x47, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1898, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1899, x0_c, x5_c, x6, x11_c, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w1900, x5_c, x9, x10, x11, x18_c, x26_c, x27_c, x32_c, x35_c, x38_c, x48_c, x50_c, x56, x61, x62_c, x67_c, x68_c, x74_c, x76, x80_c, x82, x84, x93_c);
and (w1901, x0, x3, x10, x13, x14, x15, x16_c, x22_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1902, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x61_c, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1903, x2_c, x3_c, x5_c, x6_c, x7_c, x8_c, x10, x11, x12, x15, x16, x17, x22_c, x25, x28_c, x29_c, x31, x33, x38_c, x39, x42_c, x45, x46_c, x47, x50_c, x51, x54_c, x55, x56, x58, x60, x61, x64, x65, x66, x70_c, x71_c, x72_c, x75_c, x78, x81, x82_c, x84_c, x85, x88, x89_c, x92_c, x93, x95_c, x96_c, x97, x98, x99);
and (w1904, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92_c, x94_c, x95_c, x97_c, x98_c, x99);
and (w1905, x49, x94_c, x95, x96, x97_c);
and (w1906, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x64_c, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w1907, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1908, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1909, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1910, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88_c, x93_c, x97_c);
and (w1911, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91_c, x93_c, x95_c, x96, x98, x99);
and (w1912, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1913, x5, x10, x16, x21_c, x34_c, x35, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w1914, x3_c, x5, x6, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1915, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79, x80_c, x82_c);
and (w1916, x0, x1, x2_c, x4_c, x5, x6_c, x8, x9, x10_c, x11, x12_c, x14, x15, x17_c, x18_c, x20_c, x21_c, x22, x23, x24_c, x25, x27, x28, x30, x32, x33, x34_c, x35, x37_c, x38, x40, x41, x42, x43_c, x44_c, x45, x46_c, x47_c, x48, x49, x50, x51, x52, x53_c, x54, x55_c, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64, x66_c, x67_c, x69, x70, x71, x74_c, x75_c, x76, x79, x80, x81_c, x83_c, x86, x87_c, x89_c, x90_c, x92, x93, x94, x95_c, x97, x98_c, x99_c);
and (w1917, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1918, x5_c, x9, x27, x61_c, x76, x77, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1919, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1920, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1921, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x62_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1922, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16, x17_c, x18_c, x19_c, x20, x21, x22_c, x23_c, x24_c, x25, x26_c, x27_c, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x35, x36_c, x38, x39_c, x41, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x54, x55_c, x56_c, x57_c, x58_c, x59, x60, x61, x62, x63_c, x64_c, x65, x66_c, x68, x69, x70_c, x71, x72, x73_c, x74_c, x77, x79_c, x80, x81_c, x82, x83_c, x86_c, x87_c, x88_c, x89, x90, x91_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w1923, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89, x93_c, x97_c);
and (w1924, x0_c, x1, x2, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1925, x12_c, x15_c, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1926, x5_c, x9, x26, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1927, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1928, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1929, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x69_c, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w1930, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x54_c, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1931, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1932, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1933, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1934, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x22, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1935, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w1936, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1937, x0_c, x5, x23_c, x28_c, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1938, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84, x93_c, x97_c);
and (w1939, x0_c, x1_c, x3, x4_c, x5, x6_c, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1940, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x93_c, x95_c, x96, x98, x99);
and (w1941, x1, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11, x12, x13_c, x15_c, x16_c, x17, x18_c, x19, x20, x21, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31, x32_c, x33_c, x34_c, x35_c, x36, x37_c, x38_c, x39, x40, x41, x42, x44_c, x45, x46, x47, x48_c, x49, x50, x51_c, x52, x53, x54, x55, x56, x57_c, x58, x59_c, x65_c, x67_c, x68_c, x69, x70_c, x71, x72, x73_c, x74, x76_c, x77, x78_c, x79, x80_c, x81_c, x82, x83_c, x85_c, x86_c, x87, x88_c, x89_c, x90, x91_c, x92, x93_c, x95, x97, x98);
and (w1942, x18_c, x24, x25_c, x26, x28_c, x30, x31_c, x34_c, x36, x42_c, x48_c, x51_c, x53, x56_c, x59_c, x79_c, x80, x81_c, x83, x92_c, x94, x95, x99_c);
and (w1943, x32_c, x51, x60);
and (w1944, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x64, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w1945, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56_c, x73_c, x76, x85, x89, x93, x97_c);
and (w1946, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81_c, x90_c, x93_c, x97_c);
and (w1947, x3, x4, x5_c, x6, x7, x8, x10_c, x14_c, x16_c, x17, x18, x24_c, x25_c, x27, x28, x29, x31, x34, x36, x37, x38_c, x41_c, x42_c, x45, x47, x48, x49, x53_c, x54, x57_c, x58_c, x59_c, x60_c, x63_c, x64_c, x66_c, x67_c, x68_c, x69, x74_c, x76_c, x78, x81, x82_c, x85_c, x91_c, x92, x96_c, x98_c, x99_c);
and (w1948, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x75, x77, x82, x83, x93_c, x97_c);
and (w1949, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x79, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1950, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87_c);
and (w1951, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w1952, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44_c, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1953, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x95, x97_c);
and (w1954, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x75_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1955, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x43_c, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1956, x6, x17_c, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1957, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x42_c, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w1958, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1959, x0, x1, x2_c, x4_c, x5, x6_c, x7, x8, x9, x11_c, x12, x13_c, x14_c, x15, x16_c, x17, x19, x20, x21_c, x22_c, x23, x25, x26, x27_c, x28, x29_c, x30, x31, x33, x34, x35, x37_c, x38, x40, x41_c, x42, x45_c, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62_c, x64_c, x65_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75_c, x76, x77, x81, x82_c, x83, x84, x85_c, x86, x88_c, x90_c, x91_c, x93, x94, x95_c, x96, x97_c, x98_c);
and (w1960, x0, x1, x4_c, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1961, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1962, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76_c, x77, x82, x83, x93_c, x97_c);
and (w1963, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1964, x0, x1_c, x2_c, x4, x5, x6_c, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w1965, x0, x4_c, x15_c, x18_c, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1966, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41_c, x71_c);
and (w1967, x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6, x7, x8, x9, x10, x11, x12_c, x13_c, x14, x15_c, x16, x17_c, x18_c, x19, x20, x21_c, x22, x23, x24_c, x25, x26, x27, x28, x29_c, x30_c, x31, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39, x40, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47_c, x48, x49, x50, x51, x52_c, x53_c, x54, x55_c, x56, x57, x58_c, x59_c, x60, x61, x62_c, x63, x64, x65, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80_c, x81_c, x82_c, x83_c, x84_c, x85, x86_c, x87, x88_c, x89, x90, x91, x92, x93_c, x94, x95, x96_c, x97_c, x98_c, x99_c);
and (w1968, x0_c, x2_c, x3, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1969, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w1970, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
assign w1971 = x13_c;
and (w1972, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78_c, x83_c);
and (w1973, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x48, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w1974, x0, x1_c, x2_c, x4, x5, x6, x8, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w1975, x0, x2, x5_c, x6, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1976, x1, x3_c, x7, x12_c, x13, x14, x15_c, x20_c, x21_c, x22, x25_c, x26, x28, x33_c, x37, x46, x48_c, x50, x55, x62, x64, x65, x72, x75, x81, x84, x90_c, x93, x95_c);
and (w1977, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w1978, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1979, x13_c, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1980, x2, x14_c, x15_c, x17_c, x21_c, x22, x25_c, x32_c, x37, x46, x47, x49, x55_c, x56, x57, x60, x71, x72, x80, x83, x86, x88_c, x90, x95_c);
and (w1981, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w1982, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1983, x12_c, x21_c, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1984, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w1985, x5_c, x9, x10, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1986, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94, x95, x96_c);
and (w1987, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x73, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w1988, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w1989, x3_c, x5_c, x6_c, x7, x8_c, x9, x14_c, x15, x17_c, x18, x19_c, x21_c, x22, x23, x25, x26_c, x27_c, x28, x30_c, x31_c, x32, x33, x35_c, x36, x38_c, x39_c, x41_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48, x49_c, x50, x52, x53_c, x54, x55, x56, x57_c, x58_c, x59, x60_c, x62, x63_c, x64_c, x65_c, x67_c, x68, x69, x70, x71, x72_c, x73_c, x74_c, x76, x77, x78, x79_c, x80, x81_c, x82, x83_c, x84, x86, x87_c, x88_c, x89_c, x90_c, x92, x94, x95, x96, x97, x98);
and (w1990, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x75_c, x77, x82, x83, x93_c, x97);
and (w1991, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w1992, x12_c, x32, x33, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w1993, x6, x16, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w1994, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x60, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w1995, x0, x1, x2_c, x3, x5_c, x7, x9, x10, x11_c, x13_c, x17, x18, x19_c, x20_c, x21, x25_c, x27, x28_c, x29, x32, x33_c, x35_c, x36, x42_c, x43_c, x44, x46, x48_c, x49_c, x51_c, x52_c, x54_c, x56, x58_c, x60, x63_c, x64, x66_c, x68, x70_c, x74, x75, x77_c, x80_c, x81_c, x82, x83, x86, x88, x89, x91_c, x92, x95, x97);
and (w1996, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w1997, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x94_c, x95, x96_c, x98, x99_c);
and (w1998, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x89, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w1999, x0, x2, x3, x5, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2000, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x45_c, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2001, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61_c, x71_c);
and (w2002, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2003, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2004, x0, x3, x4_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2005, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x46, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w2006, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2007, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68, x75, x84_c, x85_c, x97_c);
and (w2008, x4, x38_c, x41, x78_c, x85);
and (w2009, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x64, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2010, x0, x1_c, x2_c, x3_c, x4, x5_c, x6, x7_c, x8, x9_c, x10, x11, x12_c, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x20, x21, x22_c, x23_c, x24, x25, x26_c, x27, x28, x29, x30, x31, x32, x33_c, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43_c, x44, x45, x46_c, x47_c, x48_c, x49, x50, x51, x52_c, x53, x54, x55_c, x56, x57_c, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75, x76_c, x77, x78, x79, x80_c, x81, x82_c, x83, x84, x85_c, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93_c, x94, x95, x96, x97, x98_c, x99);
and (w2011, x0, x3, x10, x13, x14_c, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2012, x5_c, x9, x27, x61_c, x62_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2013, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x58, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2014, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x90_c, x93_c, x96_c, x97, x99_c);
and (w2015, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2016, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2017, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x86_c, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2018, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x75_c, x77, x82, x83, x88, x93_c, x95_c);
and (w2019, x0, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w2020, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x52, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2021, x0, x3, x10, x13, x14, x15, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2022, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2023, x0, x2_c, x3_c, x4_c, x5, x6_c, x7, x8, x9, x10, x11_c, x13, x14_c, x15, x16, x17, x19_c, x20, x21_c, x22, x23_c, x24, x25, x26_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35_c, x36, x37_c, x38, x39, x40_c, x43_c, x44, x45_c, x46_c, x47_c, x48_c, x49_c, x50, x51_c, x52, x53, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62_c, x63, x64, x65_c, x67, x68, x69_c, x70, x71, x73, x74_c, x75, x77_c, x78, x79_c, x80_c, x81_c, x82, x83, x84_c, x85_c, x87, x88, x89_c, x90_c, x91, x92, x93_c, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w2024, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x61, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2025, x2_c, x5_c, x6_c, x7, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2026, x3, x13, x24, x27_c, x29, x31_c, x32, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2027, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x32, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2028, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x53, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2029, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2030, x1_c, x2, x3, x5_c, x6, x8_c, x9, x11_c, x12_c, x13_c, x17, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35_c, x36, x37, x38, x40_c, x42_c, x47_c, x48, x49, x54_c, x56_c, x59, x63, x64_c, x67, x68, x69_c, x70_c, x73_c, x74_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84, x86_c, x87_c, x90, x92, x94, x95, x96_c, x97, x98);
and (w2031, x0, x6, x9, x11_c, x14, x15_c, x21, x22, x24, x31, x33_c, x35_c, x41, x44_c, x49, x53, x60, x62, x65_c, x66_c, x79, x83, x91_c, x93_c, x94_c);
and (w2032, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w2033, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2034, x1, x2, x3, x4_c, x5, x7_c, x9_c, x10_c, x11_c, x12_c, x14_c, x16_c, x17_c, x18_c, x19, x20, x21_c, x22, x24_c, x25, x30, x31_c, x32, x37_c, x38_c, x40, x41_c, x42_c, x43, x44_c, x45, x48, x49_c, x50, x52, x53_c, x55, x57_c, x58_c, x59, x61, x65, x69_c, x70, x71, x72_c, x73, x74_c, x75_c, x76, x77, x78, x79_c, x81_c, x82, x86, x87, x88_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c);
and (w2035, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x27_c, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2036, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x42, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w2037, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2038, x12_c, x40, x82, x90_c, x95_c, x96_c, x98, x99_c);
and (w2039, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2040, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2041, x0, x3, x4, x8_c, x9, x10_c, x12, x16, x17, x20_c, x23_c, x24, x25, x26, x27_c, x28, x29_c, x30_c, x33, x35_c, x36, x38_c, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x50_c, x51_c, x52, x53, x54, x55_c, x56, x58_c, x59_c, x63_c, x65, x66, x67_c, x68_c, x70_c, x73_c, x76, x78, x79, x80_c, x82_c, x84, x85, x89, x90, x92_c, x93_c, x94_c, x96_c, x98);
and (w2042, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x51_c, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2043, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2044, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x68_c, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2045, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44, x71_c);
and (w2046, x9_c, x17_c, x24, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2047, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x75, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2048, x9_c, x17_c, x23, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2049, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19_c, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2050, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2051, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50_c, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2052, x5_c, x9, x27, x42_c, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2053, x0, x7, x9_c, x12, x13_c, x16_c, x20, x23, x35, x57_c, x58, x70, x75_c, x95);
and (w2054, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w2055, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2056, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79, x80_c, x82, x83);
and (w2057, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2058, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x77, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2059, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x80, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2060, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x88, x90_c, x91, x92, x95, x97_c);
and (w2061, x2, x4_c, x6, x7, x8_c, x9, x11, x12, x13, x14, x15, x16, x17, x19_c, x20, x21_c, x23_c, x24, x25, x26, x27_c, x28, x29, x31_c, x32_c, x35_c, x36_c, x38_c, x41_c, x42_c, x44, x45, x46_c, x47_c, x50_c, x51, x52_c, x53, x54, x55_c, x56_c, x59, x61, x62, x65_c, x66, x67_c, x68, x69, x71_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x81_c, x82, x83, x84, x85_c, x86, x87_c, x88, x90, x92_c, x93_c, x95_c, x97_c, x98_c);
and (w2062, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2063, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2064, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x85_c, x86_c, x87, x88_c, x89, x90, x92, x93, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2065, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x44_c, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2066, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84_c, x88, x89, x90_c, x92_c, x93, x95_c);
and (w2067, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2068, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2069, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88_c, x90_c, x93_c, x97_c);
and (w2070, x14, x17, x22, x25_c, x33, x39_c, x45, x63, x69, x77_c, x83_c, x84_c, x97_c);
and (w2071, x1, x3, x5_c, x49, x50_c, x64_c, x66_c, x70_c, x73, x79, x89, x92_c, x96);
and (w2072, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x68, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2073, x5_c, x9, x27, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2074, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2075, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x95, x96_c, x98, x99_c);
and (w2076, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x35_c, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2077, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2078, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2079, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2080, x0_c, x2_c, x8, x9_c, x10_c, x11, x13, x14_c, x15, x16, x17_c, x18_c, x19, x21, x25, x27_c, x28_c, x29_c, x30, x31_c, x34_c, x35, x36_c, x37_c, x38, x39, x41, x42_c, x43_c, x44, x45_c, x46_c, x49, x50, x51_c, x52, x53, x54_c, x55_c, x56_c, x58, x60_c, x63, x64_c, x65, x66, x67, x69, x71_c, x72, x73_c, x74, x75, x77_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x86_c, x89, x90_c, x92, x93_c, x98);
and (w2081, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x84_c, x85_c, x97, x98, x99_c);
and (w2082, x0_c, x4_c, x5_c, x6_c, x7, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2083, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x50, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2084, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2085, x1, x2, x3, x6_c, x7_c, x8_c, x10, x11, x12, x14_c, x15, x19_c, x20, x21_c, x22, x26, x28_c, x29, x30, x31, x35_c, x36_c, x38, x39, x43_c, x45, x47, x48_c, x52_c, x56, x60_c, x61, x64, x66_c, x69_c, x72_c, x73, x75, x76, x77, x79, x80, x81_c, x83, x93, x95_c, x97_c, x99);
and (w2086, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2087, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2088, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2089, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2090, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2091, x0_c, x3_c, x4, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w2092, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2093, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2094, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74_c, x79, x90_c, x93_c, x97_c);
and (w2095, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w2096, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2097, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x43, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2098, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2099, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x40_c, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2100, x0_c, x1, x2, x3_c, x4, x5, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2101, x0_c, x2_c, x4_c, x7, x8, x14_c, x15_c, x17, x21_c, x23_c, x28_c, x29, x31, x36_c, x40_c, x41, x46, x48, x52, x53, x57_c, x59_c, x62, x63_c, x64_c, x67, x68_c, x74_c, x77_c, x78_c, x79_c, x81, x82_c, x83_c, x84_c, x88_c, x96_c);
and (w2102, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x51_c, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2103, x4, x6, x7_c, x8, x10_c, x16_c, x29, x35, x36, x38_c, x45, x51, x53, x54_c, x56, x57, x66, x69, x72_c, x73_c, x74, x76, x78, x79, x82_c, x83, x84_c, x85, x86_c, x88, x92_c);
and (w2104, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2105, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x94, x95_c, x96, x97_c);
and (w2106, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2107, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x93_c, x95_c, x96, x98, x99);
and (w2108, x0, x1_c, x2, x3, x4, x5, x6, x7, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23, x24, x25, x26_c, x27_c, x28, x29, x30_c, x31, x32, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40, x41, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x63_c, x64, x65, x66, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75_c, x76_c, x78, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95_c, x96, x97, x98, x99);
and (w2109, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18_c, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2110, x49, x92_c, x94_c, x95_c, x96, x97_c);
and (w2111, x1, x3, x5_c, x6_c, x8_c, x9, x10_c, x11_c, x12, x13, x16_c, x18_c, x19, x21_c, x22, x23, x25_c, x26_c, x27_c, x28_c, x30, x31, x34, x36_c, x37_c, x38_c, x39, x40_c, x41_c, x42, x43_c, x44, x47_c, x48, x50_c, x51, x55_c, x57, x58_c, x59_c, x60, x63, x64, x65_c, x66, x69, x70_c, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x80, x81_c, x82, x83_c, x84_c, x85, x88_c, x89, x90, x91_c, x92_c, x94, x95, x96, x97_c, x98);
and (w2112, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x18, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2113, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85, x89, x93, x97_c);
and (w2114, x2_c, x11, x29_c, x53_c, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2115, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x76, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2116, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x75_c, x77, x82, x83_c, x88_c, x93_c, x95_c);
and (w2117, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2118, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2119, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34_c, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2120, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91_c, x95, x99);
and (w2121, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91, x92_c, x93_c, x95_c, x96, x98, x99);
and (w2122, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2123, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70_c, x82, x90_c, x96, x98, x99_c);
and (w2124, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59_c, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2125, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x32_c, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2126, x0_c, x1_c, x2, x3_c, x8_c, x10, x11_c, x12, x16, x18_c, x20, x21, x22, x23, x26, x27, x30, x31, x32_c, x33, x34, x39_c, x44_c, x47, x55_c, x58, x60, x62, x66_c, x67, x69_c, x74, x75_c, x77_c, x82_c, x85, x93_c, x95_c, x98, x99_c);
and (w2127, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x71_c, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2128, x3_c, x4, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2129, x1_c, x2, x3_c, x4, x5, x6_c, x7_c, x8, x9_c, x11, x12_c, x13, x14_c, x15, x16_c, x17_c, x18_c, x19_c, x20, x21, x23, x24_c, x25_c, x26, x27, x28, x29, x30_c, x31_c, x32, x33_c, x34, x35_c, x36_c, x38, x39_c, x40_c, x41_c, x42, x43, x44_c, x45, x46_c, x47, x48, x49, x50, x51, x52_c, x53, x54, x55_c, x56_c, x57_c, x58_c, x60, x61, x62, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x73, x74, x75, x76_c, x77_c, x78, x79, x80_c, x81_c, x82, x83, x84, x85_c, x86, x87, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97, x98_c, x99_c);
and (w2130, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2131, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2132, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x91_c, x92, x95, x97_c);
and (w2133, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96_c, x97, x98_c);
and (w2134, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x85_c, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w2135, x73, x81, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2136, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54_c, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2137, x0, x1, x2_c, x3, x4, x5_c, x6_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w2138, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x91_c, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2139, x0, x4_c, x13, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2140, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2141, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70, x71_c);
and (w2142, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x66_c, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2143, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2144, x0_c, x3_c, x4_c, x6_c, x12_c, x40, x82, x90_c, x96, x98, x99_c);
and (w2145, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2146, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w2147, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2148, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x77_c, x79_c, x82, x93, x97_c);
and (w2149, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x90, x91, x92, x95, x97_c);
and (w2150, x1, x2_c, x3, x6_c, x7, x8_c, x9, x11, x12_c, x14_c, x15_c, x17_c, x18, x19_c, x20, x24_c, x27, x29_c, x31_c, x35_c, x40, x41, x42, x44, x46_c, x48_c, x49_c, x51, x52_c, x56_c, x58, x60_c, x62, x63, x68_c, x69, x71_c, x73, x74_c, x75_c, x76_c, x79_c, x81, x82_c, x84_c, x85_c, x88_c, x89_c, x93_c, x94_c, x95_c, x96_c, x97, x99_c);
and (w2151, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x65_c, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2152, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2153, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2154, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2155, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x44, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2156, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2157, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2158, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x84, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2159, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91);
and (w2160, x12_c, x40, x80, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2161, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w2162, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2163, x0_c, x1, x2, x3, x7, x8, x9_c, x10_c, x11, x12, x13_c, x14_c, x15, x17, x18, x20, x21_c, x22, x23_c, x24_c, x25, x26_c, x27, x29_c, x30_c, x31_c, x32, x33_c, x35, x36, x37_c, x39, x40_c, x41_c, x42_c, x43, x44, x47_c, x48_c, x49, x50, x52, x53, x54, x56_c, x57, x58_c, x59, x60, x61, x63_c, x64_c, x65, x66_c, x68_c, x69, x70, x72_c, x73, x74_c, x76, x77_c, x79, x80, x81, x85, x86, x87, x88, x89, x91_c, x92, x95_c, x96, x97, x99);
and (w2164, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x28_c, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2165, x4_c, x5_c, x7_c, x8, x9_c, x10, x83_c);
and (w2166, x0, x2, x7, x15_c, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2167, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w2168, x0_c, x1_c, x4, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x18, x19, x20_c, x21, x23_c, x26_c, x27, x30_c, x31, x32_c, x33, x34, x35, x38, x42, x48, x49_c, x50_c, x51_c, x53, x56_c, x61_c, x62_c, x66, x67, x68_c, x69_c, x72, x75_c, x76_c, x77_c, x79_c, x80, x81_c, x83_c, x84, x85_c, x86_c, x87, x89_c, x91_c, x93, x94, x95, x96, x98);
and (w2169, x0_c, x1, x2_c, x7_c, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14_c, x15, x16, x18, x19, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26, x27, x29, x30, x31_c, x34, x35, x36, x37, x38_c, x40_c, x41, x42, x44_c, x45_c, x46_c, x48, x49, x50_c, x51_c, x53, x54, x55, x56_c, x57, x58_c, x59, x60, x62_c, x64_c, x65, x66, x67_c, x68_c, x70, x71, x72_c, x73_c, x74, x75_c, x76_c, x77, x80_c, x81, x83_c, x84, x85, x86, x87, x90, x91, x92_c, x93_c, x94, x95_c, x98, x99_c);
and (w2170, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2171, x3, x13, x19_c, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2172, x0, x1, x2, x4, x9, x10_c, x11_c, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2173, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2174, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x83, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2175, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36_c, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2176, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91, x92, x93_c, x94, x96_c, x97_c);
and (w2177, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2178, x0, x2, x3, x6_c, x10_c, x11, x13_c, x15, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2179, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x96_c, x97, x98, x99_c);
and (w2180, x7, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2181, x0_c, x5, x23_c, x25, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2182, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2183, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2184, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x93_c, x95_c, x96, x98, x99);
and (w2185, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2186, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2187, x44_c, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2188, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2189, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2190, x12_c, x32, x70, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2191, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x87_c, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2192, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x63, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2193, x11, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2194, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x49, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2195, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2196, x1, x2_c, x4, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2197, x0_c, x3, x4_c, x5_c, x7, x8_c, x9_c, x10_c, x12, x17, x20, x22, x24, x26_c, x27_c, x28_c, x33, x38_c, x39_c, x42_c, x43, x44, x45_c, x46_c, x47_c, x48, x49_c, x51, x52, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61, x63_c, x64, x65, x70, x73_c, x74, x77_c, x78, x79, x80, x83_c, x85_c, x86, x88, x89_c, x93, x94_c, x95, x97_c, x98_c, x99);
and (w2198, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2199, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2200, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x68_c, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2201, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25, x40, x82, x90_c, x96, x98, x99_c);
and (w2202, x0_c, x2_c, x4, x5, x7_c, x9_c, x13_c, x14, x16_c, x18, x21, x23_c, x24_c, x25_c, x26, x27_c, x31, x34, x35, x37, x44, x45, x49, x50_c, x51, x52_c, x54, x59_c, x60, x61_c, x64, x65, x68, x70, x71, x73_c, x74, x78_c, x80_c, x81_c, x82, x86, x88, x92_c, x93_c, x94_c, x95_c, x97, x99_c);
and (w2203, x1, x2_c, x6, x7_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2204, x13_c, x14_c, x17, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w2205, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2206, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2207, x0_c, x1, x4_c, x5_c, x6, x8, x10_c, x12, x14, x16_c, x18_c, x19, x20_c, x21, x22_c, x23_c, x25, x27_c, x29_c, x30, x33, x34, x36_c, x38_c, x39, x44, x45, x47, x49_c, x51, x52, x54_c, x56, x59, x61, x62_c, x63, x66, x67, x68, x69_c, x70_c, x75_c, x77, x78, x79_c, x80_c, x83_c, x84, x86, x87, x89, x90, x91, x92, x93_c, x94, x95, x96_c, x97, x99);
and (w2208, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w2209, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2210, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90_c, x93_c, x97_c);
and (w2211, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56_c, x83_c);
and (w2212, x11_c, x14_c, x16, x18_c, x24_c, x31_c, x38, x43_c, x45, x47_c, x48_c, x52_c, x62, x65, x70_c, x80, x83_c, x86_c, x87_c, x89_c, x95, x99_c);
and (w2213, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x83_c, x93_c, x97_c);
and (w2214, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x53, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2215, x0_c, x5, x6, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2216, x1, x2, x3_c, x6_c, x9_c, x10, x11_c, x14_c, x17, x18_c, x20, x22_c, x24_c, x28, x29_c, x32_c, x36_c, x38, x39, x42_c, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x52_c, x56, x59, x60_c, x61, x62_c, x65_c, x66_c, x67_c, x68, x73_c, x77, x78_c, x79_c, x85_c, x86, x87, x88, x91, x92, x93_c, x96, x97_c, x98, x99_c);
and (w2217, x0, x3, x10, x13, x14, x15, x16_c, x22, x23, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w2218, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2219, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x72_c, x79, x90_c, x93_c, x97_c);
and (w2220, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2221, x5_c, x9, x27, x61_c, x67_c, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2222, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x65_c, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2223, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x19, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2224, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2225, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w2226, x5_c, x9, x27, x61_c, x76, x86, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2227, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2228, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2229, x0, x1_c, x2, x5_c, x7, x8, x9, x10_c, x12, x13_c, x14_c, x15_c, x16_c, x17_c, x18, x20, x22, x23_c, x24, x25, x26, x27, x28_c, x29, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x38, x39, x40, x41_c, x42, x43_c, x45, x46_c, x47_c, x48_c, x50_c, x51_c, x52, x53, x56, x57_c, x58_c, x59_c, x61_c, x62, x64, x65_c, x66, x67_c, x68_c, x69, x70_c, x71, x72, x73_c, x74, x77, x78, x79_c, x80, x81_c, x82, x84_c, x85, x86, x87, x88, x89, x91_c, x92_c, x93, x94, x95, x96_c, x97_c, x99_c);
and (w2230, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2231, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x77_c, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2232, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2233, x28, x34, x37, x38_c, x40_c, x44, x46_c, x47, x53_c, x67_c, x69, x73, x76_c, x78, x80_c, x81, x91, x94, x99);
and (w2234, x0, x1_c, x7, x9, x10_c, x12, x13_c, x14, x16, x19, x20, x21, x22_c, x24, x25_c, x26, x29, x30, x34_c, x35_c, x36_c, x37, x38_c, x41, x43, x48, x50_c, x52, x53_c, x54_c, x55, x56_c, x57_c, x58_c, x61_c, x65_c, x66, x67, x68_c, x69, x70, x72, x73_c, x75_c, x77_c, x78, x79, x83_c, x84, x86_c, x87_c, x89_c, x90_c, x92_c, x93, x94, x95, x98_c);
and (w2235, x4_c, x10, x15_c, x22_c, x23, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w2236, x1, x3, x4_c, x5, x7, x8, x9_c, x10_c, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2237, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2238, x5_c, x9, x12_c, x13, x14, x25_c, x32_c, x35_c, x47, x48, x50, x58_c, x63_c, x67_c, x75, x80, x86_c, x93, x94, x95_c, x96);
and (w2239, x0_c, x1_c, x2_c, x4, x5_c, x6_c, x7, x8, x9, x10_c, x11, x12, x13_c, x15_c, x16_c, x19_c, x21_c, x23, x24, x27, x28_c, x30_c, x32, x33_c, x34, x36_c, x37, x38, x39, x41, x42, x45_c, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x54, x55, x57, x58_c, x59_c, x60, x61_c, x62, x63_c, x64_c, x65, x66, x67, x68, x69_c, x70, x73, x75_c, x76_c, x77_c, x78, x79_c, x80, x81_c, x82, x84_c, x85, x86, x87, x89_c, x90, x91_c, x93_c, x94, x95_c, x97, x98, x99_c);
and (w2240, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x70_c, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2241, x8_c, x14_c, x23, x26, x38, x51_c, x62_c, x70, x77_c, x92_c, x99_c);
and (w2242, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2243, x0, x4_c, x15_c, x22_c, x25_c, x30, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2244, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x43_c, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2245, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55, x73_c, x76, x85, x89, x93, x97_c);
and (w2246, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2247, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x79, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2248, x0_c, x3, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2249, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2250, x9_c, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2251, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2252, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38, x40, x82, x90_c, x96, x98, x99_c);
and (w2253, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2254, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2255, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x84_c, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w2256, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x70, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2257, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x20_c, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2258, x1, x2, x5_c, x7, x9_c, x12, x13_c, x15_c, x23_c, x26, x28, x30, x38, x40, x45_c, x52_c, x53_c, x55, x59_c, x67, x68, x69_c, x73, x74, x80, x83, x84_c, x89, x90, x92_c);
and (w2259, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2260, x12, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2261, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2262, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x89_c, x93, x97_c, x98_c, x99_c);
and (w2263, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
assign w2264 = x29;
and (w2265, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x80_c, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2266, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x45, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2267, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2268, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2269, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18_c, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2270, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2271, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2272, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51_c, x82, x90_c, x96, x98, x99_c);
and (w2273, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x83_c, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2274, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74, x82, x90_c, x96, x98, x99_c);
and (w2275, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x83, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2276, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2277, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47, x83_c);
and (w2278, x0, x2_c, x3_c, x4_c, x5, x7_c, x9, x11_c, x12, x14_c, x15_c, x18, x21_c, x22, x28, x30_c, x31, x32, x34, x35_c, x37, x38, x39_c, x43, x47_c, x49_c, x50, x51_c, x52, x55_c, x59, x60, x63, x66, x68_c, x72_c, x75_c, x76_c, x78, x82_c, x84_c, x88_c, x89, x90_c, x91, x92, x93_c, x95_c, x96);
and (w2279, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x97_c, x98, x99_c);
and (w2280, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2281, x0_c, x5, x23_c, x30_c, x31, x32_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2282, x0_c, x1, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2283, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2284, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7_c, x8, x9_c, x10, x11, x12, x13_c, x14_c, x15, x16_c, x17_c, x18_c, x19, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x34, x35, x36, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55_c, x56_c, x57_c, x58, x59_c, x60, x61_c, x62, x63_c, x65_c, x66_c, x67, x69_c, x70_c, x71_c, x72, x73_c, x75_c, x76_c, x77, x78, x79, x80, x82_c, x83_c, x84_c, x85, x86_c, x87_c, x88, x89_c, x90, x91, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w2285, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x56_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2286, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2287, x0, x3, x10, x13, x14, x15, x16_c, x22, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2288, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x34_c, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2289, x3, x12, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2290, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2291, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2292, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2293, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x61_c, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2294, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x92_c, x95, x97_c);
and (w2295, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2296, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x63, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2297, x8, x12, x18, x24_c, x27, x35_c, x39_c, x47_c, x51, x58, x62, x79, x80_c, x83);
and (w2298, x2, x4_c, x6, x8_c, x11_c, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2299, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2300, x49, x66, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2301, x0, x1, x6_c, x7, x10_c, x12_c, x14_c, x15, x17_c, x18_c, x21, x24_c, x25, x28, x30, x32, x36_c, x39, x41_c, x44, x48, x51_c, x54, x55, x56, x58_c, x59, x60_c, x61, x62, x64_c, x65, x66_c, x68_c, x69_c, x70, x73_c, x74, x77, x79, x81_c, x82, x83, x87, x88, x89_c, x92_c, x93_c, x94, x95_c, x97_c, x98, x99);
and (w2302, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x24, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w2303, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x10_c, x12, x13, x14, x15_c, x16_c, x17_c, x18_c, x19, x20_c, x21, x22, x23_c, x24, x25, x26_c, x27_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36_c, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49_c, x50, x51_c, x52, x53, x54, x55, x56, x57, x58_c, x59, x60, x61_c, x63, x64_c, x66_c, x68, x69, x70_c, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x79, x81_c, x82, x84, x85, x86, x87, x88, x89_c, x90_c, x91, x92_c, x93, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w2304, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2305, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x39_c, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2306, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2307, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x60_c, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2308, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2309, x2_c, x11, x29_c, x31, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2310, x0_c, x1, x2_c, x4, x5, x9_c, x10_c, x12_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19, x20_c, x21_c, x22_c, x24, x25_c, x26_c, x28, x29, x30_c, x32, x33_c, x34, x35, x36_c, x37_c, x38, x39, x40, x42, x43, x44, x45_c, x46, x47, x48_c, x50_c, x51_c, x52, x53_c, x55_c, x56, x57, x59, x60_c, x62, x63_c, x64, x66, x67_c, x68, x69_c, x71, x72_c, x73, x74_c, x75_c, x76_c, x78_c, x81_c, x83_c, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93, x95_c, x96, x97_c, x98_c, x99);
and (w2311, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2312, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2313, x0_c, x1, x4_c, x5_c, x8, x9_c, x10, x11_c, x13_c, x14, x15_c, x16_c, x17, x18, x19_c, x21_c, x22, x24, x25_c, x28_c, x29_c, x31_c, x32_c, x33, x34, x35, x36, x37, x38_c, x39, x40, x41, x43_c, x47_c, x49, x50, x51, x52_c, x54_c, x55_c, x56_c, x57, x58, x61_c, x62, x63, x64_c, x65, x67_c, x70_c, x73, x74_c, x75, x76_c, x77, x78, x79, x81, x83, x84, x86_c, x88, x89_c, x90_c, x92_c, x93, x98_c, x99_c);
and (w2314, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2315, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85_c);
and (w2316, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2317, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2318, x13_c, x14_c, x37_c, x39_c, x45_c, x51_c, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2319, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x83_c, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2320, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x58, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2321, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x87_c, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2322, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2323, x36, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2324, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2325, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2326, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86);
and (w2327, x2_c, x19, x24_c, x26, x36, x46_c, x55_c, x92_c, x95_c, x98);
and (w2328, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58, x83_c);
and (w2329, x31_c, x36, x38_c, x47, x63, x67_c, x69_c, x75_c, x89);
and (w2330, x12_c, x40, x70_c, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2331, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x28_c, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2332, x1, x6, x14, x19_c, x26_c, x33_c, x48, x53, x59_c, x70, x76, x78_c, x83, x95_c);
and (w2333, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96, x97_c);
and (w2334, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2335, x12_c, x40, x82, x90_c, x98_c, x99_c);
and (w2336, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2337, x23, x39, x55_c, x64, x65, x70, x74);
and (w2338, x2, x4_c, x5, x6, x7_c, x9_c, x13, x14, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2339, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2340, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88, x90_c, x93_c, x94, x95, x96, x97, x98, x99);
and (w2341, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x30_c, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2342, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x45_c, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2343, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2344, x0_c, x1_c, x2_c, x9_c, x10_c, x12, x13, x21_c, x25, x26_c, x27_c, x34_c, x39_c, x45_c, x48, x53, x55, x56_c, x60, x64, x70_c, x72, x74_c, x76_c, x78_c, x79_c, x80, x82_c, x84_c, x85_c, x88, x89, x90, x94_c, x95, x98_c, x99);
and (w2345, x0_c, x1_c, x3, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2346, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x57, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2347, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2348, x1, x2_c, x3, x4_c, x7, x8_c, x9, x13_c, x14_c, x15, x17, x18_c, x24_c, x26, x31_c, x33, x35, x36_c, x38, x39, x40, x41_c, x42_c, x43, x44_c, x50_c, x52, x56_c, x58_c, x62_c, x65_c, x67, x70, x72_c, x73_c, x75, x76_c, x77_c, x79_c, x80, x81_c, x82, x84_c, x85_c, x86, x88, x92_c, x94_c, x96_c, x97_c, x99_c);
and (w2349, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2350, x8, x21_c, x25_c, x27_c, x34, x39_c, x41_c, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2351, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2352, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2353, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2354, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x67_c, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2355, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x93_c, x96, x97_c);
and (w2356, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2357, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2358, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2359, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x65, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2360, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2361, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x84_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2362, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2363, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x47_c, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2364, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2365, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x75, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2366, x62_c, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2367, x0, x1, x2, x3, x4, x5, x7_c, x8, x9_c, x11, x13_c, x15, x16_c, x18, x19_c, x20_c, x24_c, x25, x26_c, x27_c, x29_c, x30, x31_c, x33_c, x34, x35, x36_c, x37, x38, x39, x41, x43, x45, x47_c, x48_c, x53_c, x55, x57, x58_c, x59_c, x61, x62, x64_c, x65_c, x66_c, x69, x71, x72_c, x74_c, x76_c, x77, x78_c, x81_c, x82_c, x83_c, x84_c, x85_c, x87_c, x88, x89_c, x91, x95_c, x96, x97_c, x99_c);
and (w2368, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x70_c, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2369, x8, x21_c, x25_c, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2370, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x25, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2371, x0, x5, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2372, x6_c, x7, x8_c, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2373, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x77, x82, x83, x93_c, x97_c);
and (w2374, x2, x5, x6_c, x7_c, x8, x12, x16, x17, x19_c, x21_c, x25_c, x27_c, x29_c, x30_c, x35, x36, x38_c, x39_c, x42_c, x47_c, x50, x51_c, x52_c, x53, x58_c, x59, x65_c, x70_c, x72_c, x73, x76_c, x78, x79, x81_c, x82_c, x83, x85_c, x90_c, x91_c, x93_c, x94, x95, x97, x99);
and (w2375, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2376, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x33, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2377, x0, x1_c, x2_c, x4, x5, x6, x8, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2378, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2379, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x88_c, x90, x93_c, x95_c, x96, x98, x99);
and (w2380, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2381, x0_c, x1, x3_c, x4, x6_c, x8, x9_c, x11_c, x13_c, x15_c, x17_c, x19_c, x21, x23, x24_c, x28_c, x29_c, x30_c, x31, x32_c, x33, x34, x36, x39, x41, x42_c, x47_c, x49_c, x50_c, x54, x56_c, x58, x59_c, x60, x61_c, x62_c, x63_c, x64, x65_c, x70, x73_c, x74, x75, x77, x80, x81, x83_c, x84_c, x87, x88, x89, x91, x92_c, x93, x95_c, x97_c, x98_c);
and (w2382, x0, x2, x3, x4_c, x5, x6_c, x7, x8, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19_c, x20, x21_c, x22_c, x24_c, x25, x26, x27, x28, x30_c, x31, x32_c, x33_c, x34, x36, x37_c, x38, x40_c, x41, x42_c, x43_c, x45, x47_c, x48, x49, x50, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x57_c, x58, x59, x60_c, x61, x62, x63, x64_c, x66, x67, x69, x70_c, x71, x72_c, x74, x75, x76_c, x77_c, x78_c, x79, x80, x81, x82_c, x83_c, x84_c, x86, x87_c, x88_c, x89_c, x90, x91, x92_c, x93_c, x94_c, x95_c, x96, x97, x98, x99);
and (w2383, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2384, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x61_c, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2385, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w2386, x0_c, x3, x5, x7_c, x8, x9_c, x10, x11, x12, x13_c, x14_c, x15_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x25, x26, x28, x29_c, x30, x31_c, x32, x33, x34_c, x35_c, x36, x37_c, x39, x40_c, x42, x43, x44, x45_c, x46, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61, x62, x63, x64_c, x65, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x73, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83_c, x84, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92, x93_c, x94_c, x95_c, x96_c, x98_c, x99);
and (w2387, x2, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w2388, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x52, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2389, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2390, x1_c, x2, x3_c, x4, x5_c, x6_c, x8_c, x9_c, x10_c, x11_c, x14, x16_c, x18, x20, x22_c, x23, x24, x25, x28_c, x30_c, x31, x32_c, x33, x37, x39, x40, x41_c, x43, x45_c, x46_c, x47, x49, x50, x51, x52, x53, x55, x56, x57_c, x58_c, x59_c, x60, x62, x63_c, x64_c, x66_c, x67, x68_c, x70_c, x71, x72, x74, x75_c, x77, x78, x80, x81, x82, x83, x84, x85, x86_c, x87_c, x89, x90_c, x91, x93_c, x94_c, x95, x97_c);
and (w2391, x0, x1_c, x4, x5, x6_c, x7, x8, x9, x11, x12_c, x13_c, x15_c, x16, x18_c, x20, x21, x22, x23, x24, x25, x26_c, x29_c, x30, x31_c, x32, x33_c, x35_c, x36_c, x37_c, x38, x39, x40, x41_c, x44_c, x45, x46, x47, x49, x50_c, x51, x52_c, x53_c, x54_c, x55_c, x56, x57_c, x58, x59, x60, x61, x63, x64, x65, x66, x68_c, x69, x70, x71, x74_c, x76_c, x78, x80_c, x81_c, x82, x83_c, x85, x90_c, x92_c, x93, x94_c, x96_c, x98);
and (w2392, x0_c, x1, x3, x4_c, x5, x6, x7_c, x8_c, x10, x11_c, x12_c, x14, x15_c, x16_c, x17, x18, x20_c, x21_c, x22_c, x23_c, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31_c, x32, x33_c, x34_c, x36_c, x38, x39_c, x40_c, x41, x43, x44_c, x46, x47_c, x48_c, x50, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x57, x58, x60, x61_c, x62, x63_c, x64_c, x65, x66, x67_c, x70_c, x71, x72, x73_c, x75, x76_c, x79_c, x80_c, x81_c, x82, x83_c, x84_c, x85, x86, x87_c, x88, x92_c, x93, x94_c, x95_c, x96, x97_c, x98, x99);
and (w2393, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x56_c, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2394, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2395, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x91, x92_c, x93, x94, x95, x97_c, x99_c);
and (w2396, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2397, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2398, x0, x1, x2_c, x4_c, x6_c, x7, x8_c, x12, x13, x15, x16_c, x21_c, x25_c, x27_c, x28, x30, x31, x33_c, x34_c, x35, x37, x38_c, x39, x40, x42, x43, x44_c, x47_c, x49_c, x52, x54_c, x55, x56, x58_c, x59, x61_c, x62_c, x64, x66, x67, x68, x69, x70_c, x74, x75, x76, x77, x80, x81, x84, x85_c, x86_c, x90, x91_c, x94, x95, x97, x98);
and (w2399, x23, x46_c, x51_c, x58);
and (w2400, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2401, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x92_c, x93_c, x94, x95, x96, x99);
and (w2402, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2403, x21_c, x35_c, x41, x57, x59_c, x62_c, x73_c, x85_c, x91);
and (w2404, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2405, x0_c, x1, x2_c, x3_c, x5_c, x7_c, x8_c, x11_c, x12, x14_c, x15, x16_c, x17_c, x20_c, x23_c, x24_c, x25, x26_c, x28_c, x29, x32, x34, x35, x36, x37_c, x38, x40_c, x42, x43, x44_c, x45, x47_c, x48_c, x49, x50_c, x51_c, x52, x56_c, x57_c, x58, x61, x62, x68_c, x69_c, x71, x74, x76, x77_c, x78_c, x79, x80_c, x81_c, x83, x84_c, x86, x87_c, x88, x89_c, x90, x92_c, x94, x95, x96_c, x97_c, x98_c, x99_c);
and (w2406, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2407, x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16_c, x19, x20, x21_c, x22, x23, x24_c, x25_c, x27, x28, x29, x30, x32, x33_c, x34, x35_c, x36, x37, x38_c, x39, x40, x41_c, x42, x43, x44_c, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52_c, x53, x54, x55_c, x56, x57_c, x58, x59_c, x60, x61_c, x62, x63_c, x64, x66_c, x67_c, x69, x70_c, x71_c, x73_c, x74, x76_c, x77_c, x78, x79, x80, x81_c, x82_c, x83, x84_c, x85_c, x86, x87, x88_c, x89_c, x90, x91, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98, x99_c);
and (w2408, x0_c, x1_c, x2_c, x3, x4_c, x5, x6, x7_c, x8_c, x9, x10_c, x11_c, x12, x13, x14, x15_c, x16, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x24, x25_c, x26_c, x28_c, x29, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38_c, x39_c, x41, x42, x43_c, x44, x45, x46, x47_c, x48, x49, x50_c, x51, x52, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x68, x69, x70, x71_c, x72_c, x73_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93, x94_c, x95, x96, x97_c, x98, x99);
and (w2409, x1_c, x2_c, x3_c, x4, x5_c, x8, x9_c, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2410, x1_c, x2_c, x4, x5_c, x9_c, x10, x11_c, x13, x15_c, x16_c, x21, x23, x24, x25_c, x26, x28_c, x31, x34, x37_c, x42, x43, x46, x47, x48_c, x49, x50, x53_c, x54, x55, x56, x57, x59_c, x61_c, x64, x65, x70, x73_c, x75, x77_c, x78_c, x80, x81_c, x83, x85, x86, x90, x91, x94, x96);
and (w2411, x4, x5, x9, x15, x19_c, x23, x29, x32_c, x33_c, x38, x40_c, x42_c, x50_c, x62_c, x63_c, x69, x70_c, x73, x74, x79_c, x81, x82_c, x86_c, x91_c, x92_c, x97_c);
and (w2412, x0_c, x2, x3_c, x8_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2413, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2414, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2415, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x87, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2416, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x61_c, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2417, x0_c, x1, x3_c, x5_c, x6, x7, x8, x9, x10, x11_c, x12_c, x14, x15_c, x16, x17_c, x18, x20_c, x21, x22, x23_c, x25, x26_c, x27, x28_c, x31_c, x32, x33, x35_c, x36_c, x37, x38_c, x39, x42, x46_c, x47_c, x49_c, x51_c, x52_c, x53_c, x54, x55, x56_c, x57, x59_c, x60_c, x62, x63_c, x64, x66, x69_c, x70_c, x71, x72_c, x75, x77_c, x80_c, x81_c, x82_c, x84, x85_c, x86_c, x87_c, x89, x90, x91_c, x93, x94, x99_c);
and (w2418, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98_c);
and (w2419, x2_c, x11, x24, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2420, x0, x2, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2421, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2422, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x38_c, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2423, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x64_c, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2424, x0_c, x2_c, x3_c, x4_c, x6, x7, x8, x9_c, x10_c, x11, x12_c, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x24, x25, x26_c, x27, x28, x29, x30_c, x31_c, x32, x33, x34, x35, x36_c, x38, x40_c, x41, x42, x43, x44, x45_c, x46_c, x47, x48_c, x49, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57, x58_c, x59, x60, x61, x62, x63_c, x64_c, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x74, x75, x76_c, x77_c, x79, x80, x81_c, x82_c, x83, x84, x86_c, x88_c, x89, x90, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w2425, x0, x7, x8, x12, x14, x28, x33_c, x34, x40_c, x41, x55, x58_c, x61_c, x62, x68_c, x72, x77, x80_c, x82, x84_c, x87, x92_c, x97_c);
and (w2426, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x98_c, x99);
and (w2427, x0, x5_c, x6, x10_c, x11_c, x15, x17, x18, x19_c, x20_c, x21_c, x22, x27_c, x29_c, x30_c, x32, x33_c, x34, x36_c, x37, x42, x45_c, x46_c, x48_c, x50_c, x54, x59, x60_c, x61_c, x62, x69, x70, x73, x74_c, x78_c, x80, x81, x83_c, x85_c, x86, x90, x91_c, x92, x95_c, x97_c, x99);
and (w2428, x2_c, x3, x4, x5_c, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2429, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x77_c, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2430, x3, x6, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2431, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2432, x2, x5_c, x6, x8_c, x11_c, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2433, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2434, x0_c, x5, x23_c, x30_c, x31, x32, x38, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2435, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2436, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x77_c, x82, x83, x93_c, x97_c);
and (w2437, x3, x5_c, x7_c, x8_c, x11_c, x14_c, x15_c, x16_c, x17, x18_c, x20, x21, x22_c, x24_c, x29_c, x30_c, x31_c, x32, x33, x34_c, x39, x41, x52_c, x54, x55, x56_c, x57_c, x58, x63_c, x64, x68_c, x69_c, x79_c, x82_c, x83_c, x84_c, x86_c, x88, x89, x90_c, x95, x96, x97_c);
and (w2438, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x10, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2439, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x52_c, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2440, x1_c, x2_c, x3_c, x6_c, x8, x9, x11_c, x12, x14, x15, x18, x20, x21, x23, x26_c, x27, x29, x31_c, x32, x34_c, x36, x39_c, x40_c, x41, x44, x45, x47_c, x48, x49_c, x52, x53_c, x54, x55_c, x57_c, x58_c, x63_c, x66, x68_c, x69_c, x70, x72_c, x74_c, x75, x77, x78, x83_c, x84_c, x86_c, x87, x89, x91, x92, x93_c, x94, x96_c, x98);
and (w2441, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2442, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x72, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2443, x0_c, x4, x13_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2444, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2445, x0_c, x2, x4_c, x7, x10, x15, x16_c, x20_c, x22_c, x23_c, x29, x30, x31_c, x37_c, x41, x44_c, x48_c, x51_c, x52, x54_c, x55, x56, x57, x61_c, x62, x65, x70, x73, x74, x75_c, x78, x79_c, x81, x85, x88, x91_c, x93, x99_c);
and (w2446, x1_c, x4, x5_c, x6_c, x7_c, x10_c, x14_c, x16, x17_c, x19_c, x20, x22_c, x25, x26_c, x27_c, x28, x30_c, x32, x33, x34_c, x35_c, x37, x38_c, x41, x43_c, x44, x48_c, x51, x52, x53, x55, x56, x58, x59_c, x60_c, x66, x70, x71_c, x73, x78_c, x79_c, x81_c, x82_c, x83, x84, x86, x88, x89, x92, x93_c, x94_c, x96_c, x97_c, x99);
and (w2447, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2448, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2449, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x81, x84, x85, x95, x99);
and (w2450, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x40, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2451, x4, x83_c);
and (w2452, x5_c, x9, x27, x31_c, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2453, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2454, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2455, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2456, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x84, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2457, x1, x2, x3, x4_c, x8_c, x9, x13_c, x14, x17, x18, x19_c, x20_c, x21, x24, x26, x28, x29_c, x30_c, x31_c, x32_c, x33, x34, x37, x38_c, x40, x41, x43_c, x47, x48_c, x49, x51, x52_c, x54_c, x55, x56_c, x59_c, x60, x61_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x70, x72, x73, x75, x77, x78, x79, x80_c, x81, x82_c, x84_c, x87, x89_c, x90_c, x91, x92, x93_c, x94_c, x95, x98, x99);
and (w2458, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2459, x0_c, x1_c, x2_c, x4_c, x5_c, x6, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2460, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66_c, x83_c);
and (w2461, x0_c, x1_c, x2_c, x3, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2462, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2463, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2464, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x75_c, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2465, x0, x50_c, x51, x53, x67_c, x79, x81);
and (w2466, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2467, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2468, x5, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2469, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x80_c, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2470, x2_c, x11, x29_c, x35_c, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2471, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91, x92, x93_c, x94_c, x95, x97, x98, x99);
and (w2472, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x90_c, x92_c, x94, x97, x99_c);
and (w2473, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x69_c, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2474, x0_c, x1, x2, x4_c, x5, x6, x7, x8, x9_c, x10, x12, x13_c, x14, x15, x17_c, x18, x19_c, x20, x21_c, x24, x25, x26, x27_c, x28, x30_c, x32, x33, x34, x35_c, x36, x39_c, x42, x43, x45_c, x46_c, x47_c, x48_c, x50_c, x51_c, x53_c, x54_c, x56_c, x57, x58, x59, x60, x61_c, x62_c, x65_c, x66_c, x68, x69, x70, x71_c, x73_c, x74, x75_c, x76_c, x77, x79, x80_c, x81, x82_c, x83, x84, x85, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x94_c, x95_c, x96_c, x97, x98, x99);
and (w2475, x48_c, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2476, x2_c, x11, x29_c, x93, x95_c, x96, x98, x99);
and (w2477, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x49, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2478, x0, x1_c, x2, x3, x4_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12_c, x16, x18, x19, x20_c, x22_c, x25, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36, x37, x38_c, x39, x40, x42_c, x44, x45_c, x46, x47, x48, x49, x50, x52_c, x54, x55_c, x58_c, x59_c, x60_c, x61_c, x62_c, x64, x65_c, x66, x67, x68_c, x71_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81_c, x83_c, x84_c, x86, x88, x89_c, x91, x93, x95, x96, x97, x98_c, x99);
and (w2479, x8, x21_c, x23, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2480, x3, x11_c, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2481, x2_c, x11, x29_c, x33, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2482, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x39, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2483, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x30_c, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2484, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x47, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2485, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x64_c, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2486, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61_c, x82, x90_c, x96, x98, x99_c);
and (w2487, x12_c, x32, x61_c, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2488, x1, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2489, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87_c, x88, x89_c, x90_c, x92, x95, x97_c);
and (w2490, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x89, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2491, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2492, x1_c, x2, x4_c, x7, x9_c, x10, x11_c, x12_c, x15, x17_c, x18, x19_c, x20, x22, x24_c, x25, x26_c, x27, x28_c, x29, x30, x31, x32, x34_c, x36_c, x39_c, x40_c, x44, x46_c, x47, x49_c, x50_c, x51, x52_c, x53_c, x55_c, x56, x58_c, x59, x60, x63, x65_c, x67_c, x68_c, x69, x70, x71, x73_c, x74, x78_c, x79_c, x80, x86, x87, x88, x89, x90_c, x93, x94, x96, x97, x98_c, x99);
and (w2493, x12_c, x32, x67_c, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2494, x2, x3_c, x4_c, x5, x6, x7_c, x8, x11_c, x12_c, x15_c, x17_c, x18, x20_c, x21_c, x23, x24, x25, x26, x28_c, x29_c, x30_c, x31_c, x33, x34_c, x35_c, x39_c, x40_c, x41, x42, x43, x44, x46_c, x48_c, x50_c, x51, x52, x53_c, x54_c, x55_c, x56, x57, x58, x60_c, x61, x62, x63, x64, x65_c, x66_c, x67_c, x68, x69, x70, x71, x72_c, x73, x74_c, x75, x76, x77, x78, x79_c, x80_c, x82, x83_c, x84, x85_c, x86, x88, x89_c, x90, x91, x92_c, x94_c, x95, x96_c, x97, x98);
and (w2495, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x62, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2496, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2497, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x95, x97, x98, x99_c);
and (w2498, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2499, x1, x3_c, x4_c, x7_c, x9_c, x11, x19, x23_c, x27, x28, x29_c, x36, x37, x40, x42_c, x46_c, x48_c, x49, x50, x52, x55, x57, x58_c, x62_c, x64_c, x65, x67_c, x69, x70_c, x74, x76, x80_c, x85, x87_c, x90_c);
and (w2500, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2501, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2502, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61_c, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2503, x0, x1_c, x2, x3_c, x4_c, x5_c, x6_c, x7, x8, x9, x10_c, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17, x18, x19_c, x20, x21_c, x22, x23, x24, x25, x26, x27, x28, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36, x37, x38_c, x39_c, x40, x41, x42, x43_c, x44, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51, x52, x53, x54, x55_c, x56_c, x57, x58, x59_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68, x69_c, x70, x71_c, x72, x73_c, x74_c, x75_c, x76, x77, x78_c, x79, x80, x81, x82, x83, x84_c, x85, x86_c, x87, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98, x99);
and (w2504, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x49, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2505, x0, x4_c, x5, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2506, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w2507, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94, x95, x96, x97, x99_c);
and (w2508, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x49, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2509, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x91_c, x93_c, x94_c, x95_c, x96, x97_c, x99_c);
and (w2510, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2511, x54, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2512, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2513, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2514, x10_c, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w2515, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96_c, x97_c);
and (w2516, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x60_c, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2517, x2_c, x11, x29_c, x84_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2518, x3_c, x5, x6, x7_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2519, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x71_c, x72_c, x79, x90_c, x93_c, x97_c);
and (w2520, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x37, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2521, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2522, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2523, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2524, x13_c, x34, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w2525, x2, x5_c, x6, x9_c, x12_c, x16_c, x24, x28, x31, x33, x36_c, x39, x40, x41, x42_c, x45_c, x49, x50, x55_c, x58_c, x59, x62, x64, x66, x70, x71, x73, x80_c, x83, x88_c, x92_c, x95);
and (w2526, x18, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2527, x0_c, x1_c, x2, x3_c, x6, x8, x9, x10, x11, x12, x13, x15, x16, x18_c, x20_c, x21, x22_c, x23, x26, x28, x31_c, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x40, x43_c, x44, x45_c, x49_c, x52, x53_c, x55, x57, x58, x60, x61, x63_c, x66, x68_c, x70, x71, x74, x75, x76_c, x77, x79_c, x81, x82, x84, x85, x86_c, x88, x89_c, x91_c, x92, x93_c, x94, x95_c, x96, x98);
and (w2528, x2_c, x5, x23, x24, x39, x60, x66, x68_c, x70, x84_c);
and (w2529, x0, x1, x2_c, x3_c, x4_c, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2530, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55_c, x82, x90_c, x96, x98, x99_c);
and (w2531, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2532, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2533, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x23, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2534, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x68, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2535, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x19_c, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2536, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2537, x0_c, x1_c, x3, x4_c, x5_c, x6_c, x7_c, x8, x9_c, x11, x12_c, x13_c, x14, x15_c, x18, x20, x21_c, x22, x24, x26, x27, x30, x37_c, x38, x39, x40_c, x41, x42_c, x43, x46, x47, x50_c, x52_c, x55, x58, x61_c, x63_c, x64_c, x67, x69, x71, x74, x76, x78_c, x80_c, x81_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91, x92, x94_c, x96, x98, x99_c);
and (w2538, x0, x2_c, x3, x4_c, x5_c, x8_c, x10, x11, x15_c, x18, x29, x33, x40, x41_c, x47_c, x51, x52_c, x53_c, x56_c, x57, x61, x63_c, x64, x67, x69, x70_c, x73_c, x83, x84, x86_c, x87_c, x88_c, x90, x93_c, x94, x95, x97_c, x98, x99);
and (w2539, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x78_c, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2540, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92, x93_c, x95, x97_c);
and (w2541, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2542, x20_c, x21, x35, x40, x54_c, x70_c, x74_c, x90);
and (w2543, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17, x40, x82, x90_c, x96, x98, x99_c);
and (w2544, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2545, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x66, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2546, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x46_c, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2547, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2548, x49, x79, x90_c, x93_c, x97_c);
and (w2549, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x74, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2550, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53_c, x73_c, x76, x85, x89, x93, x97_c);
and (w2551, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79, x82, x83, x93_c, x97_c);
and (w2552, x3_c, x4, x5, x6_c, x8_c, x10_c, x12, x14, x15_c, x17_c, x19_c, x20, x21, x24, x29_c, x32_c, x33_c, x34, x36, x40_c, x48_c, x50_c, x55_c, x56, x60, x61_c, x62, x66, x68, x72_c, x73, x76, x78_c, x79_c, x84_c, x87, x90, x92_c);
and (w2553, x12_c, x23_c, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2554, x11, x12_c, x15, x17_c, x23_c, x26, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2555, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2556, x5_c, x9, x27, x41, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2557, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92, x93_c, x95_c, x96, x98, x99);
and (w2558, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2559, x8_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2560, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12, x13_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2561, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2562, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2563, x12_c, x13_c, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2564, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81, x82, x83, x93_c, x97_c);
and (w2565, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x67, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2566, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2567, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2568, x0_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2569, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2570, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2571, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89, x90_c, x92, x94_c, x96_c, x97, x98, x99_c);
and (w2572, x11, x12_c, x15_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2573, x5_c, x9, x27, x61_c, x74_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2574, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2575, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2576, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x39, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2577, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2578, x14, x15, x20_c, x31_c, x36_c, x42_c, x48, x59_c, x63, x64, x67_c, x70, x73_c, x74_c, x88);
and (w2579, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w2580, x8_c, x12_c, x14, x15, x18_c, x19, x23_c, x24_c, x26, x30, x32, x35, x36_c, x41_c, x47_c, x56_c, x76_c, x77_c, x78_c, x82, x90, x91_c, x98, x99);
and (w2581, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x11_c, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2582, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x57_c, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2583, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x97);
and (w2584, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83, x84_c, x85_c, x97_c);
and (w2585, x0, x3, x53_c, x59_c, x77, x82_c, x91);
and (w2586, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2587, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2588, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2589, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2590, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2591, x2_c, x4_c, x8, x9, x11, x12_c, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2592, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34_c, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2593, x0_c, x1_c, x3_c, x4_c, x5_c, x6, x7_c, x8, x9_c, x11_c, x12_c, x13_c, x15_c, x16, x17_c, x18_c, x20, x23, x24_c, x25, x26, x27_c, x28, x29, x30, x33, x34, x36, x37, x38_c, x43_c, x45_c, x46_c, x47, x49_c, x50, x51, x52_c, x54_c, x55_c, x56_c, x58, x60_c, x61, x62_c, x63_c, x64_c, x65, x66, x67, x68, x69, x70, x71, x73, x74, x79_c, x82, x84, x85, x86, x88_c, x89, x91, x93_c, x94, x96_c, x97, x98_c);
and (w2594, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2595, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x8_c, x9, x11, x12, x13_c, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x23_c, x24_c, x25_c, x27, x28, x29_c, x30, x31, x32, x33_c, x34, x35, x37, x38_c, x40, x41, x42_c, x43, x45, x47, x48_c, x49, x50_c, x51, x52, x53, x54, x55_c, x56_c, x58, x59_c, x61, x62, x63, x64, x65, x67_c, x68, x69_c, x70_c, x71, x72, x73_c, x75, x76_c, x77, x78, x79_c, x80, x81, x82_c, x83, x84_c, x85, x86, x87, x89, x91, x93, x94, x95_c, x96, x97, x98_c);
and (w2596, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2597, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x67, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2598, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2599, x0_c, x1, x2_c, x3_c, x5, x7_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16_c, x17_c, x18, x19, x20, x21, x22_c, x23, x24, x25, x26, x27_c, x28_c, x29, x31_c, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39, x40_c, x41, x42, x43, x44_c, x45, x46, x47_c, x49_c, x50, x51_c, x52_c, x53, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x67, x68_c, x69_c, x70_c, x71_c, x72_c, x73, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83, x84_c, x86, x87, x88, x89_c, x90_c, x91, x92_c, x93, x94, x95, x96_c, x97, x98, x99_c);
and (w2600, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2601, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x12, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2602, x0, x1, x2, x4, x7, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2603, x0_c, x2_c, x4_c, x7_c, x8_c, x9, x11, x12, x16, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2604, x0_c, x6_c, x9, x11_c, x19, x23_c, x26, x32, x35_c, x45_c, x48, x55, x57, x58_c, x61, x67_c, x69_c, x71, x75, x77, x80, x84_c, x85_c, x87_c, x91_c, x96_c, x97_c, x98);
and (w2605, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2606, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2607, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2608, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2609, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x70_c, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2610, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2611, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x55_c, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2612, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x93_c, x96, x97_c, x98, x99_c);
and (w2613, x12_c, x17_c, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2614, x29_c, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2615, x11, x12_c, x15, x17_c, x18_c, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2616, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2617, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2618, x1_c, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2619, x1, x2_c, x3, x4, x5, x6, x7_c, x8_c, x9_c, x11, x13_c, x14, x15, x16_c, x17, x19_c, x20, x21, x22_c, x23, x24, x26, x27_c, x29_c, x30_c, x31_c, x32_c, x33_c, x38_c, x40_c, x41_c, x43_c, x45, x47, x48_c, x49_c, x50, x52_c, x53_c, x54, x55_c, x60, x61_c, x63, x64, x67, x69_c, x70, x71, x73, x74, x75_c, x77, x78_c, x80_c, x81_c, x82, x83_c, x84_c, x85_c, x88_c, x89_c, x90, x91_c, x92_c, x93, x99);
and (w2620, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x64, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2621, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x15, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2622, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2623, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2624, x1_c, x2, x3_c, x4, x11_c, x12, x14, x15, x16, x18_c, x20, x21_c, x22_c, x24, x26_c, x27_c, x29, x30_c, x32_c, x33_c, x34_c, x35, x36, x37_c, x40, x43, x44, x47, x50_c, x52_c, x53_c, x54_c, x55_c, x56_c, x58, x59_c, x60, x63, x69, x70, x73_c, x76, x77_c, x82_c, x83_c, x84, x88, x89_c, x90, x92, x95, x97_c, x98_c);
and (w2625, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x40_c, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2626, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2627, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x90, x96, x98, x99_c);
and (w2628, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2629, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w2630, x12_c, x32, x39, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2631, x5_c, x6, x10_c, x11_c, x19_c, x20_c, x21, x23, x24, x29, x32_c, x34_c, x35, x36_c, x37, x38_c, x39_c, x44, x49_c, x53_c, x55_c, x57, x58, x59, x60, x61_c, x64, x67_c, x68_c, x70_c, x72, x74, x79, x80_c, x81_c, x83, x85, x86, x87_c, x90, x92_c, x96, x98, x99);
and (w2632, x6, x17_c, x20_c, x24_c, x25_c, x27, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w2633, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x81, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2634, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w2635, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x92, x96, x97_c);
and (w2636, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x37_c, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2637, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2638, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2639, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53_c, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2640, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89, x95, x99);
and (w2641, x0_c, x1, x3, x5, x6, x7, x9, x10_c, x13, x15_c, x17_c, x21_c, x24_c, x26_c, x28, x30, x31, x33_c, x36_c, x41, x45_c, x46_c, x47_c, x54, x56, x61_c, x64, x66_c, x67_c, x75, x78_c, x85, x86, x87_c, x88, x89_c, x94_c, x96, x97_c);
and (w2642, x0, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2643, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2644, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2645, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2646, x49, x71_c, x72_c, x79, x90_c, x93_c, x97_c);
and (w2647, x0_c, x3_c, x4_c, x6, x7_c, x10, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2648, x0, x1, x2, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2649, x3, x13, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2650, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
assign w2651 = x52_c;
and (w2652, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x59, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2653, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x96_c, x97_c, x98, x99_c);
and (w2654, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x87_c, x89, x90_c, x91_c, x93, x94_c, x96, x97);
and (w2655, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91, x92, x93_c, x94_c, x95, x96, x97, x99);
and (w2656, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2657, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79, x80_c, x82, x83_c, x84_c, x91_c, x92_c);
and (w2658, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x87, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2659, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2660, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27_c, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2661, x0, x1, x2, x3, x5, x9, x10, x12_c, x13_c, x14, x15, x17_c, x18_c, x21_c, x22_c, x24_c, x25, x26_c, x29, x30_c, x31_c, x32, x33, x36, x37_c, x38_c, x39, x41_c, x42_c, x43, x44_c, x45_c, x48_c, x49_c, x53, x54, x58, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69, x70, x71_c, x72, x74, x75_c, x76, x78_c, x79, x80, x81_c, x82, x83_c, x85, x87, x88_c, x89, x90_c, x91_c, x92_c, x93, x94_c, x95, x98_c);
and (w2662, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91, x92_c, x93_c, x97_c);
and (w2663, x1_c, x2, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x12, x13, x14, x15_c, x16, x17, x18_c, x20, x21, x22, x23, x25, x26_c, x28, x30, x31_c, x32_c, x34_c, x35_c, x36_c, x37_c, x38_c, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48_c, x49, x51, x52, x53_c, x54_c, x55, x56_c, x59, x61, x62, x63, x65, x66_c, x67_c, x68, x69_c, x70_c, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x81, x82, x83_c, x84, x85, x86_c, x87_c, x88, x89, x91_c, x92_c, x93, x94, x95, x96_c, x97, x98_c, x99);
and (w2664, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2665, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2666, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57_c, x83_c);
and (w2667, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2668, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2669, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2670, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x71_c, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2671, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2672, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2673, x0_c, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w2674, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2675, x11_c, x15, x23_c, x71_c);
and (w2676, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x25_c, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2677, x39_c, x54, x55, x58_c, x62, x71, x81_c, x94);
and (w2678, x12_c, x32, x90_c, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2679, x49, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2680, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2681, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x65, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2682, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2683, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30_c, x40, x82, x90_c, x96, x98, x99_c);
and (w2684, x0, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11_c, x12, x13_c, x14, x15, x16_c, x17_c, x18, x19_c, x20_c, x22, x23_c, x24_c, x25_c, x26_c, x27_c, x28, x29, x30_c, x31, x33_c, x34_c, x35_c, x36_c, x37_c, x38_c, x39_c, x40, x41_c, x42, x43_c, x44_c, x45, x46_c, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x55, x56_c, x57_c, x58, x59_c, x60, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x72_c, x73, x74, x75_c, x76, x77, x78_c, x79, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88_c, x89, x90, x91, x92_c, x93, x96_c, x97, x98, x99);
and (w2685, x18_c, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2686, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2687, x3_c, x12_c, x16_c, x20, x44_c, x52, x66, x69_c, x92_c);
and (w2688, x6, x17_c, x20_c, x24, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w2689, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x89, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2690, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2691, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2692, x43_c, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2693, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91_c, x93_c, x95_c, x96, x98, x99);
and (w2694, x0, x2, x5_c, x6_c, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2695, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2696, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2697, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x88, x90_c, x91, x92, x95, x97_c);
and (w2698, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x65, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2699, x13_c, x14_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2700, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2701, x0, x1, x2, x4, x9_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2702, x4_c, x6_c, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w2703, x2, x11_c, x31, x35, x42_c, x81, x97_c, x99_c);
and (w2704, x13_c, x14, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2705, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2706, x2_c, x9, x12_c, x14, x17_c, x20, x23_c, x28_c, x41_c, x46, x53_c, x63, x64_c, x75, x79_c, x80_c, x82_c, x84, x92, x93_c);
and (w2707, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x98, x99_c);
and (w2708, x49, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2709, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x87, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2710, x0, x4, x6_c, x7_c, x9_c, x12_c, x14_c, x16, x19_c, x22, x24_c, x25, x26_c, x27, x31, x35, x37_c, x38, x41_c, x42, x43_c, x44, x45_c, x46, x47, x49_c, x53, x55, x56_c, x61, x64_c, x65, x70_c, x71_c, x72, x74, x76_c, x77, x79_c, x82, x84, x87, x89_c, x90_c, x93_c, x94, x95_c, x96_c, x97_c);
and (w2711, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x30, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2712, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w2713, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2714, x0, x1_c, x2, x3_c, x4, x5, x6_c, x7_c, x9, x10, x12_c, x13_c, x14, x15_c, x16, x19_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x40_c, x41_c, x42_c, x43, x45_c, x47, x48_c, x51_c, x52, x53_c, x54_c, x56, x58_c, x59, x60_c, x61, x62, x63, x66, x67_c, x69, x74, x75, x76_c, x77_c, x78, x79, x80_c, x81, x83_c, x84, x88, x89, x92, x94_c, x95_c, x96_c, x97_c, x99_c);
and (w2715, x0, x1, x2_c, x6_c, x7_c, x8_c, x10, x12, x14_c, x15_c, x16_c, x17_c, x19, x20_c, x22, x24, x25_c, x27, x31_c, x32_c, x33, x34_c, x37_c, x38, x39_c, x40_c, x41, x42, x43, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51_c, x53, x54, x55, x56_c, x57, x58, x60_c, x61, x62_c, x64_c, x66, x67_c, x70_c, x71_c, x72, x73, x75_c, x76_c, x80_c, x81_c, x83_c, x85_c, x92, x93_c, x99_c);
and (w2716, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x87, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2717, x0_c, x1_c, x2, x3_c, x4_c, x5, x6_c, x8_c, x9_c, x10_c, x11, x12_c, x13_c, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29, x30_c, x31_c, x32, x33_c, x34_c, x36_c, x37_c, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53_c, x54, x55_c, x56_c, x57_c, x58, x59_c, x60, x61_c, x62, x63_c, x64_c, x65_c, x66_c, x67, x68, x69_c, x70_c, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81, x82, x83_c, x84_c, x85, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94, x95_c, x96_c, x97, x98_c, x99);
and (w2718, x4_c, x20_c, x25_c, x33_c, x34, x41_c, x43_c, x46_c, x50, x54, x66, x69, x72_c, x77_c, x80, x82, x86);
and (w2719, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2720, x0_c, x16, x38, x53_c, x84, x99);
and (w2721, x2_c, x4_c, x5, x9, x10, x11, x13, x15, x16, x20, x21, x22_c, x23_c, x25, x26_c, x27, x28_c, x31_c, x33, x36_c, x40, x44_c, x47, x52_c, x62, x63, x65_c, x68, x69, x72_c, x73, x74, x76, x78, x81, x83, x84, x85, x87_c, x88, x89, x94, x95);
and (w2722, x73, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2723, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2724, x2_c, x3, x4, x6_c, x11_c, x13_c, x14, x15_c, x18_c, x19_c, x20_c, x22_c, x23, x25, x27, x29_c, x30, x32_c, x33_c, x34_c, x39_c, x40, x43, x44_c, x47_c, x49, x50_c, x52, x53, x56, x60, x62_c, x66, x67, x68_c, x72_c, x73_c, x74_c, x75, x77_c, x78, x80, x81, x82, x84_c, x85_c, x86, x87, x90, x93, x95, x96_c, x97_c);
and (w2725, x3_c, x17, x49_c);
and (w2726, x2_c, x11, x29_c, x73_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2727, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x56_c, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2728, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2729, x8, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2730, x0, x1_c, x2_c, x3, x4, x5, x6_c, x10, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2731, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x62_c, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2732, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x47, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
assign w2733 = x23_c;
and (w2734, x0_c, x1_c, x3, x4_c, x5, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2735, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2736, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87);
and (w2737, x11_c, x15_c, x16, x18_c, x23_c, x71_c);
and (w2738, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x87, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2739, x2_c, x11, x22_c, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2740, x13_c, x14_c, x23_c, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w2741, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x89, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2742, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x84_c, x85, x90_c, x96, x98, x99_c);
and (w2743, x11, x12_c, x15, x17_c, x20, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2744, x0_c, x1_c, x3, x4_c, x6, x7_c, x8, x10_c, x12, x13, x14, x18, x19, x20, x21_c, x24_c, x25, x27, x28, x29, x30, x31_c, x32_c, x34, x37, x38_c, x39, x41_c, x44, x49_c, x54_c, x56_c, x59_c, x60, x62, x63, x64_c, x65_c, x66, x67_c, x68_c, x70, x71_c, x73, x74_c, x76_c, x77, x78_c, x82, x85, x90, x91, x93, x94, x96, x97);
and (w2745, x0, x1_c, x2_c, x4, x5, x6_c, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2746, x1_c, x3, x4_c, x5, x6_c, x7, x8, x9_c, x11_c, x14, x15, x16, x17, x18, x19_c, x20_c, x22_c, x23_c, x24, x25_c, x27, x28, x29, x30, x31_c, x34_c, x35_c, x36_c, x37, x38_c, x39, x40_c, x41_c, x42, x43, x44, x46_c, x47, x49_c, x50, x51, x52_c, x53_c, x54_c, x55_c, x56_c, x58_c, x59, x60, x63, x64_c, x65_c, x66_c, x68_c, x69, x70, x71_c, x72_c, x73, x78, x79, x80_c, x81_c, x82_c, x83_c, x84_c, x85, x86, x88_c, x89, x92_c, x93_c, x94_c, x95_c, x96_c, x98_c, x99);
and (w2747, x11_c, x27, x37, x50, x51, x55_c, x57, x59, x64, x66_c, x71, x75_c, x76, x79_c, x86_c, x99_c);
and (w2748, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w2749, x0, x1, x2_c, x3_c, x6_c, x7_c, x9, x11, x12, x14, x16, x17_c, x18_c, x19_c, x20, x21_c, x22, x23, x24, x25_c, x26, x27_c, x28, x29, x30, x31_c, x32, x33, x34_c, x35_c, x36_c, x37, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52_c, x53, x54, x56_c, x57, x58_c, x59, x60, x61_c, x62, x63_c, x64, x65, x66, x67, x68, x69, x70_c, x71_c, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x84, x85, x86, x88, x89_c, x90_c, x91_c, x94, x96, x97_c, x98_c, x99_c);
and (w2750, x9_c, x17_c, x26, x27, x28_c, x29_c, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2751, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2752, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2753, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2754, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92, x93, x97_c);
and (w2755, x1, x7, x8, x10_c, x16, x20, x22_c, x29_c, x36, x39, x45, x47, x51_c, x52_c, x55, x57, x60, x61, x66_c, x72, x74, x75_c, x91_c, x98);
and (w2756, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x20, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2757, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x83_c, x93_c, x97_c);
and (w2758, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2759, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x92_c, x95, x97_c);
and (w2760, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96, x99);
and (w2761, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34, x83_c);
and (w2762, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2763, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2764, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x85, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2765, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2766, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2767, x10, x13_c, x14, x30, x33_c, x34_c, x42_c, x45, x51, x56_c, x64, x68, x71_c, x72_c, x73_c, x75_c, x77, x79, x80_c, x94);
and (w2768, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85_c, x93_c, x97_c);
and (w2769, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x28, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2770, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x89, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2771, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x35, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w2772, x0_c, x5, x23_c, x29_c, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2773, x1_c, x41, x55, x65_c, x74_c, x89, x94_c);
and (w2774, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2775, x16, x38, x55, x63, x77, x82_c, x93);
and (w2776, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x21_c, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2777, x0, x4_c, x15_c, x22_c, x25_c, x27, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2778, x2_c, x21, x62, x81_c, x98);
and (w2779, x0_c, x2_c, x3_c, x6_c, x7, x8, x9_c, x10, x11_c, x12_c, x13_c, x14, x16_c, x17, x18, x19_c, x22_c, x23_c, x24_c, x27, x28_c, x29, x31, x32_c, x33, x34, x35, x36, x38, x39, x40_c, x41_c, x42, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51_c, x54, x55, x58, x59, x60, x61_c, x63, x64, x65_c, x66_c, x67_c, x69_c, x70, x71, x72, x73_c, x74, x75_c, x77_c, x78, x79, x81_c, x82, x83_c, x84, x85_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99);
and (w2780, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2781, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w2782, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2783, x2_c, x3_c, x4, x6, x7, x8, x9_c, x10, x11, x12_c, x13, x16, x17_c, x18_c, x19_c, x21_c, x22, x24_c, x25, x26, x28_c, x29, x30, x31_c, x32, x33, x34, x35, x36_c, x38, x39, x40, x41_c, x42_c, x45_c, x46, x48, x50_c, x51_c, x54_c, x55, x56_c, x60_c, x61, x62, x63, x64_c, x65, x66, x67, x68_c, x70_c, x71, x72, x76, x77_c, x78_c, x79, x80, x81_c, x82, x83, x84_c, x85_c, x87_c, x88_c, x92, x93_c, x94, x95, x96, x98, x99);
and (w2784, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2785, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x80_c, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2786, x0_c, x2_c, x4_c, x5_c, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2787, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2788, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2789, x0, x1, x2_c, x3, x4_c, x5_c, x6_c, x9, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2790, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90_c, x93, x97_c);
and (w2791, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84, x90_c, x93_c, x97_c);
and (w2792, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2793, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x40, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2794, x13_c, x49, x64, x71, x72_c, x79, x81, x87, x90, x93_c, x97_c);
and (w2795, x2_c, x11, x29_c, x43, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2796, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2797, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2798, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40, x71_c);
and (w2799, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28_c, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2800, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79, x84_c, x85_c, x97_c);
and (w2801, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77_c, x83_c);
and (w2802, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2803, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x33, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2804, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x82_c, x83, x93_c, x97_c);
and (w2805, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x55, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w2806, x0, x1_c, x2_c, x4, x5_c, x6, x8_c, x10_c, x13, x14_c, x17_c, x18, x19, x20, x24, x25_c, x27_c, x28_c, x29, x30_c, x33_c, x34_c, x36, x37, x38, x40, x41_c, x46_c, x47, x49_c, x50_c, x52_c, x53, x54_c, x55_c, x56, x57_c, x63_c, x64, x65_c, x66, x67, x68, x70, x71, x73_c, x74_c, x75, x76_c, x77, x78_c, x79_c, x80_c, x83_c, x84, x85, x88, x89_c, x91_c, x92, x94, x95_c, x96, x97_c, x98_c, x99);
and (w2807, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2808, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2809, x0_c, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9, x10, x11, x12, x13_c, x14_c, x15_c, x16, x17, x18_c, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x43_c, x45, x46, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66, x67_c, x68, x69_c, x70_c, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79, x80, x81_c, x82_c, x83_c, x84, x85_c, x86, x87, x88_c, x89_c, x90, x91_c, x92, x93, x94_c, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w2810, x0_c, x1_c, x2, x3_c, x6, x7, x8_c, x9_c, x12_c, x13, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x23_c, x24, x25, x26, x27, x28, x30, x31_c, x32, x34, x35_c, x36_c, x37, x38_c, x39, x41_c, x42_c, x43_c, x44, x45_c, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x55_c, x56, x57_c, x58_c, x59, x61, x62_c, x63, x64_c, x65_c, x66_c, x67, x68, x69_c, x70, x71_c, x72, x73, x74, x75, x76, x77, x78, x80_c, x83_c, x84, x85_c, x86, x87_c, x88, x89_c, x90_c, x93_c, x94, x96, x97, x98_c, x99_c);
and (w2811, x2, x4, x8_c, x9, x10, x11_c, x12_c, x13, x14_c, x15_c, x16_c, x18, x20, x21_c, x24_c, x25, x29_c, x37, x40, x41_c, x42_c, x43_c, x44_c, x46_c, x49_c, x50, x52_c, x53_c, x55, x56, x58_c, x61_c, x63, x65, x68, x69, x70, x71_c, x73, x74, x76, x77, x78_c, x79, x81_c, x82_c, x83_c, x85, x86_c, x87, x89_c, x91_c, x92, x94_c, x98, x99);
and (w2812, x0, x1, x2_c, x3_c, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x31, x32, x33, x34_c, x35_c, x36, x37, x38_c, x39_c, x40_c, x42_c, x43_c, x44_c, x45_c, x48_c, x49_c, x51, x52_c, x54_c, x55, x56_c, x58, x59, x60, x61, x62_c, x63_c, x64_c, x65, x66, x67_c, x68_c, x69, x70, x71_c, x72_c, x73, x74, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x82_c, x84, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93, x94, x95_c, x96_c, x97, x98_c, x99);
and (w2813, x63, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2814, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2815, x0, x1, x3_c, x4_c, x5_c, x6_c, x7, x9_c, x10, x11, x14, x15, x16, x17, x18_c, x19, x20_c, x22_c, x23, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35, x36_c, x37_c, x38_c, x39_c, x41, x42_c, x43, x44, x45, x46_c, x47_c, x48, x49, x50_c, x52_c, x53, x54_c, x56_c, x58_c, x59, x60_c, x61, x62_c, x63, x64_c, x65, x66_c, x67, x68_c, x70, x71_c, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80_c, x81_c, x82_c, x83, x84, x85, x86, x87_c, x88, x89, x90, x91_c, x92, x93, x94_c, x95_c, x96_c, x97, x98_c, x99_c);
and (w2816, x8, x12, x18_c, x20_c, x30_c, x31, x32, x33, x34_c, x37, x41_c, x43_c, x44, x46_c, x47_c, x49_c, x52, x53, x54_c, x55_c, x57, x63_c, x64, x65, x66, x67_c, x70, x73, x76_c, x77_c, x78, x82_c, x85_c, x86_c, x87, x93_c, x97_c);
and (w2817, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x15, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2818, x2, x4_c, x5, x6, x7_c, x9_c, x11, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2819, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2820, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28_c, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2821, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x29_c, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2822, x5_c, x9, x27, x61_c, x76, x88_c, x90, x91, x92, x95, x97_c);
and (w2823, x0_c, x1, x2_c, x3_c, x4, x6, x7, x8, x9_c, x10, x11, x12, x14_c, x16_c, x17, x19, x21_c, x22_c, x24, x25_c, x26_c, x27, x28, x29_c, x30, x31_c, x33_c, x34, x35, x36, x37_c, x38, x39_c, x40, x42, x43, x44, x45_c, x46, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x57, x58, x59_c, x60_c, x62, x63, x64, x66_c, x67, x68_c, x70_c, x71, x72_c, x73, x74_c, x75_c, x77, x78, x82_c, x83, x84_c, x85_c, x86, x87, x88, x89, x91_c, x92, x94_c, x96_c, x97, x98_c, x99);
and (w2824, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x72, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2825, x11, x12_c, x15, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2826, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2827, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x97_c, x98, x99_c);
and (w2828, x13_c, x14_c, x37_c, x39_c, x42, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2829, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35_c, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2830, x11, x12_c, x15, x17_c, x22, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2831, x0, x1, x2_c, x3_c, x4, x5_c, x9_c, x10, x11_c, x12, x13_c, x14, x15, x17, x18, x19, x21, x23, x24, x25, x26, x27_c, x28_c, x32_c, x33_c, x34_c, x36_c, x38_c, x39, x40, x41_c, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x50_c, x51, x52, x55_c, x57_c, x58_c, x59_c, x63_c, x64, x65, x66_c, x69, x70_c, x75, x76_c, x77, x78_c, x83, x85, x86, x87, x88, x89, x91_c, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w2832, x0_c, x4, x8_c, x10, x12, x23_c, x27_c, x37_c, x39, x43_c, x46_c, x67_c, x69, x76, x81, x82_c, x84_c, x92, x95);
and (w2833, x0, x1, x2, x3, x5_c, x6_c, x7_c, x8_c, x9, x12_c, x13, x14, x15_c, x16, x17, x18, x20, x21, x24, x25_c, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x37, x38_c, x39_c, x40, x41, x43_c, x44_c, x45_c, x47, x48, x49_c, x52, x54_c, x57_c, x58_c, x59, x60, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68, x69, x70, x71_c, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84_c, x85_c, x88, x90, x91, x92_c, x93_c, x94, x99_c);
and (w2834, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2835, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2836, x6, x15, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2837, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x36, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2838, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2839, x27_c, x33, x88_c);
and (w2840, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2841, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2842, x0, x3, x10, x13, x14, x15, x16_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2843, x0, x1_c, x2, x3_c, x4_c, x5_c, x6, x7, x8_c, x10_c, x11, x12_c, x14_c, x15, x16, x17_c, x18, x19, x20_c, x21, x22_c, x23_c, x24_c, x25, x27, x28_c, x29, x30_c, x31_c, x32, x33_c, x34, x35_c, x36, x37, x40_c, x41, x42, x43_c, x44, x45, x46_c, x47, x48, x49_c, x50_c, x51, x52, x53_c, x54_c, x55, x56_c, x57_c, x58, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x69_c, x70, x71, x72_c, x73_c, x74_c, x76, x78, x79_c, x80, x81_c, x83, x84_c, x85_c, x86, x87, x88, x89_c, x90_c, x91_c, x92, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w2844, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2845, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x71, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2846, x0_c, x2, x6_c, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w2847, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w2848, x7, x9_c, x11, x12_c, x13_c, x17, x26, x27, x29_c, x30, x32, x36_c, x40_c, x41_c, x42, x43, x46, x47, x48_c, x49_c, x52_c, x53, x57, x58_c, x60, x61, x62, x63_c, x64_c, x65, x67, x68_c, x70, x71, x72_c, x73, x74, x77_c, x82_c, x83_c, x86_c, x87, x88, x89, x90_c, x92, x93_c, x94_c, x96, x97_c, x99);
and (w2849, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2850, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x95, x96_c, x97_c);
and (w2851, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x48, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2852, x8, x21_c, x25, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2853, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2854, x2, x4, x5_c, x6, x8_c, x10_c, x13, x16_c, x17_c, x21_c, x22_c, x23, x27, x34_c, x36_c, x38, x41_c, x42_c, x52_c, x56_c, x58, x59, x60, x61_c, x64, x65, x66, x68_c, x69_c, x71, x73, x75_c, x78_c, x83_c, x85, x86_c, x89, x90, x91, x92_c, x97_c, x98);
and (w2855, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14, x83_c);
and (w2856, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x17_c, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2857, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86, x87_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2858, x87, x96);
and (w2859, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2860, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2861, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x64, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2862, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2863, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2864, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2865, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2866, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33, x83_c);
and (w2867, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2868, x0_c, x1_c, x2_c, x4_c, x5, x6, x7_c, x9, x13, x14_c, x16_c, x17, x18, x20_c, x22_c, x23, x24_c, x25, x26_c, x28, x29_c, x31_c, x32_c, x35_c, x37, x38, x40_c, x41_c, x43_c, x47, x49, x50_c, x52_c, x53_c, x54, x55_c, x56, x58, x59_c, x60, x62, x63, x64, x66, x68, x69_c, x70, x71, x72, x74_c, x75_c, x76_c, x77_c, x78, x82, x85, x88, x89, x90_c, x91, x92_c, x93_c, x94_c, x95, x98_c, x99_c);
and (w2869, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w2870, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x28_c, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2871, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2872, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x94, x95, x96_c, x98, x99_c);
and (w2873, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2874, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x8, x10_c, x11_c, x12, x13_c, x14_c, x16, x17_c, x18, x19_c, x20, x21_c, x22_c, x23, x24, x25_c, x27, x28_c, x31, x32, x33, x34, x35_c, x36_c, x37, x38, x39_c, x40, x41_c, x43, x45_c, x46_c, x48_c, x49_c, x50_c, x51, x53_c, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62_c, x65_c, x66_c, x67_c, x70, x71, x72_c, x74, x76, x77_c, x78_c, x80_c, x81_c, x82, x83_c, x84_c, x85_c, x86, x87_c, x88_c, x89, x90, x92_c, x93_c, x97_c, x98_c, x99_c);
and (w2875, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2876, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2877, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2878, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2879, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2880, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72_c, x75, x84_c, x85_c, x97_c);
and (w2881, x8_c, x49_c, x75, x89_c);
and (w2882, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w2883, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w2884, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2885, x0_c, x1, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2886, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x35, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2887, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x49_c, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2888, x12_c, x32, x88_c, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2889, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2890, x12, x13, x14, x16_c, x19, x22, x27, x30_c, x44, x56, x71_c, x98_c);
and (w2891, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2892, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x37, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2893, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2894, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w2895, x8, x18, x20_c, x40, x66, x78, x80_c, x82_c);
and (w2896, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23_c, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2897, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x32_c, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2898, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x79_c, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2899, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2900, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42_c, x82, x90_c, x96, x98, x99_c);
and (w2901, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94, x97_c);
and (w2902, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x97);
and (w2903, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x70_c, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2904, x12_c, x29_c, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2905, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97, x98, x99);
and (w2906, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2907, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2908, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2909, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w2910, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x21, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2911, x5_c, x9, x11_c, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2912, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x54_c, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2913, x0_c, x1_c, x2_c, x3, x4_c, x5, x6_c, x7, x8, x9, x10_c, x11, x12, x13_c, x14, x15, x16, x17, x18, x19_c, x20_c, x21_c, x22, x23, x24, x25, x26, x27_c, x28, x29, x31, x32, x33, x34_c, x35_c, x36, x37_c, x38, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x46, x47_c, x49_c, x50_c, x51, x52, x53_c, x54, x55, x57, x58, x59_c, x60, x61_c, x62_c, x63, x64, x65_c, x66_c, x67, x68_c, x69, x70, x71, x72_c, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x90, x91, x92_c, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2914, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25_c, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2915, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2916, x3, x13, x18_c, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2917, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w2918, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2919, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93, x95, x97_c);
and (w2920, x20, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2921, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2922, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w2923, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x96_c, x97_c);
and (w2924, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2925, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2926, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x26_c, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2927, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x97, x99);
and (w2928, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2929, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84, x93_c, x97_c);
and (w2930, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2931, x2_c, x4_c, x6_c, x7_c, x9, x11, x12_c, x14, x16_c, x18, x20_c, x21_c, x22_c, x23_c, x24, x25, x26, x27_c, x28, x32_c, x33, x36, x37_c, x39, x41, x43, x45_c, x51, x52, x53, x54_c, x56_c, x57_c, x58_c, x61, x62, x66_c, x68_c, x69_c, x71_c, x73_c, x74_c, x75, x76, x77, x80_c, x81_c, x84, x85, x86_c, x94, x96_c, x98_c, x99_c);
and (w2932, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14_c, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2933, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x70, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2934, x0, x2_c, x5, x6, x12, x15, x20_c, x24_c, x28, x31, x33_c, x35_c, x36_c, x37, x38_c, x44_c, x46, x47_c, x50, x51_c, x52_c, x55_c, x56, x58_c, x65, x69, x72, x73, x83_c, x90_c, x92, x99);
and (w2935, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w2936, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x45_c, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2937, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95_c, x97_c, x98_c, x99_c);
and (w2938, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94, x95, x96, x97, x98_c, x99);
and (w2939, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2940, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2941, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x85_c, x86_c, x87, x88_c, x89, x90, x92, x94, x95, x96_c, x97_c, x98_c, x99_c);
and (w2942, x0_c, x1_c, x4_c, x10_c, x11_c, x16, x20_c, x25_c, x34, x35, x36, x50, x54, x55, x59_c, x64_c, x69_c, x70_c, x71, x81, x86_c, x90_c, x91, x92, x93_c, x96_c);
and (w2943, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2944, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2945, x2, x4_c, x5, x6, x7_c, x9, x11_c, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2946, x0_c, x4_c, x5_c, x6_c, x8_c, x11_c, x12_c, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2947, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x64, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2948, x0_c, x2_c, x4_c, x8, x11, x14_c, x17_c, x18_c, x19, x20_c, x22, x24_c, x25_c, x26, x27, x28, x32, x33, x35_c, x36, x39, x41_c, x45, x46, x47_c, x48_c, x49_c, x51_c, x52_c, x53, x54_c, x55, x56, x58_c, x59_c, x67_c, x68_c, x71_c, x73_c, x75_c, x76_c, x77, x78_c, x82_c, x83_c, x85, x87_c, x88_c, x89_c, x90, x93_c, x96, x97);
and (w2949, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2950, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2951, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36_c, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2952, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x56, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2953, x7, x17_c, x18, x19_c, x20_c, x23_c, x24_c, x29_c, x30, x33, x44, x48, x52, x55_c, x57_c, x58, x66, x67, x73_c, x76_c, x77_c, x79, x80_c, x85_c, x86_c, x87, x89, x95_c, x96_c, x97_c, x99);
and (w2954, x2, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2955, x12_c, x32, x44_c, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2956, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w2957, x49, x62, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2958, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2959, x7_c, x9_c, x12_c, x14_c, x15_c, x16, x18, x19_c, x20_c, x22, x23_c, x24_c, x25, x30, x31_c, x32_c, x35_c, x36_c, x38_c, x39, x40, x41_c, x44_c, x46_c, x47_c, x48, x49_c, x51_c, x61, x62_c, x63_c, x65_c, x66_c, x68, x69_c, x71, x73, x74, x75_c, x77, x78, x79, x82_c, x84_c, x85, x88, x89, x90, x91, x92_c, x94, x96, x99_c);
and (w2960, x1, x3_c, x7_c, x9, x12_c, x13_c, x14, x16, x19, x20, x23, x25, x27, x28, x31, x33_c, x35_c, x39_c, x40_c, x41, x43_c, x47, x48_c, x49_c, x50_c, x52_c, x54, x55, x56, x58, x59_c, x66, x69, x73_c, x74_c, x76, x77, x81_c, x82_c, x83_c, x86, x87_c, x88, x89, x91_c, x92, x95_c);
and (w2961, x12_c, x32, x46, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w2962, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x94, x95, x96_c, x98, x99_c);
and (w2963, x0_c, x1_c, x3, x4_c, x5, x7_c, x8_c, x10, x11_c, x13, x14, x16, x18, x19_c, x22, x23_c, x24_c, x25, x26, x27_c, x28_c, x29, x30_c, x32, x33, x34_c, x35, x36, x37_c, x38, x39, x40_c, x41, x42, x43, x45, x46, x47, x49, x51_c, x53_c, x55, x56, x57, x58, x59, x63_c, x67, x68_c, x69, x70_c, x71, x72_c, x73, x75_c, x76, x77_c, x78_c, x80, x81, x82, x83_c, x84, x85_c, x86, x87_c, x89_c, x90, x93_c, x94, x96, x97, x99);
and (w2964, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88_c);
and (w2965, x5, x10, x16, x21, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w2966, x49, x75_c, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w2967, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2968, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x78_c, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2969, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2970, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2971, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x38_c, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w2972, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w2973, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2974, x0, x1_c, x2_c, x4, x5, x6, x8_c, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2975, x0_c, x1, x2, x3_c, x4, x5_c, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2976, x73, x98_c, x99);
and (w2977, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w2978, x0, x1, x2_c, x3_c, x4, x5, x6, x7, x8, x9, x10_c, x11, x12_c, x13_c, x14_c, x15, x16_c, x17, x18_c, x19_c, x20_c, x21, x22, x23, x24_c, x25, x26, x27_c, x28, x29, x30_c, x31_c, x32_c, x33, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x44_c, x45, x46_c, x47, x48_c, x49_c, x50_c, x51_c, x52, x53, x54_c, x56, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x66, x67_c, x68, x69_c, x70_c, x71, x72, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x84, x85_c, x86, x87_c, x88_c, x89, x90, x91_c, x92, x93_c, x94_c, x95_c, x96, x97_c, x98_c, x99_c);
and (w2979, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x82_c, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2980, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49_c, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w2981, x5, x10, x16, x21_c, x34_c, x35, x41, x42, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2982, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50_c, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2983, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2984, x0_c, x3_c, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w2985, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78, x83_c);
and (w2986, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w2987, x0, x1, x2_c, x3, x4, x5_c, x9, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2988, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x40, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w2989, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2990, x2, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2991, x0_c, x5, x22, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w2992, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w2993, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x44_c, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w2994, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w2995, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w2996, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51_c, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w2997, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w2998, x0_c, x2_c, x4_c, x5_c, x6_c, x7, x8, x12, x13_c, x14, x15, x16_c, x18_c, x19_c, x22, x23, x24_c, x25, x26, x28, x30, x31, x32, x33_c, x34, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x43, x44, x46, x47_c, x50, x51_c, x52, x53_c, x55_c, x56, x57, x58_c, x60, x62, x65, x66, x67, x68, x69_c, x70, x71, x74_c, x75, x76, x77, x78, x79, x81_c, x84_c, x85_c, x86, x88, x89, x91_c, x93, x95, x96_c, x97_c, x99);
and (w2999, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x25, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3000, x13_c, x14_c, x37_c, x39_c, x45, x82, x90_c, x96, x98, x99_c);
and (w3001, x12_c, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3002, x12_c, x40, x51_c, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3003, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3004, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3005, x0, x3, x9, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3006, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3007, x12_c, x32, x42, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3008, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x65, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3009, x2_c, x3_c, x4, x5, x6_c, x8, x9_c, x11_c, x12_c, x13, x14_c, x19_c, x21_c, x24_c, x28, x30, x31, x32, x35_c, x36, x39_c, x40_c, x41_c, x42, x43, x44_c, x45_c, x46, x48, x51_c, x52_c, x53, x54, x55, x57, x60_c, x61_c, x62, x63, x65_c, x68, x69, x72_c, x73, x76, x78, x79_c, x81, x82, x84_c, x86_c, x87, x90, x94, x95, x96, x97, x98);
and (w3010, x7_c, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3011, x9_c, x17_c, x21_c, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3012, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x75, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3013, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3014, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33, x40, x82, x90_c, x96, x98, x99_c);
and (w3015, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x36, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3016, x1_c, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3017, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3018, x0, x4_c, x15_c, x16, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3019, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3020, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x52, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3021, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x93_c, x95_c);
and (w3022, x2, x3, x4, x6, x7, x8, x9_c, x12, x14, x15, x16_c, x17_c, x18, x19_c, x20_c, x21, x22_c, x24, x25, x26, x27_c, x28_c, x29_c, x30_c, x33, x35, x36, x38, x40_c, x42_c, x44_c, x45_c, x47_c, x48_c, x49_c, x50, x51_c, x55_c, x56_c, x57_c, x58, x59, x61, x62_c, x64_c, x65, x67, x68, x69, x70, x71, x72, x73, x77, x78_c, x79, x80, x81_c, x82, x84, x86_c, x88, x89_c, x90_c, x91_c, x93, x94_c, x95, x96);
and (w3023, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3024, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x86, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3025, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64, x83_c);
and (w3026, x1, x2_c, x3_c, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3027, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3028, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x66, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3029, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3030, x8, x21_c, x25_c, x27_c, x34, x38_c, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3031, x0, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3032, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x78_c, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3033, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x53_c, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3034, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3035, x0, x2, x7_c, x8_c, x11, x13, x15_c, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3036, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89, x91_c, x92_c, x94, x95);
and (w3037, x1_c, x2, x6, x11, x12_c, x13_c, x20, x21, x30_c, x32, x37, x42, x49_c, x50_c, x52, x54, x55_c, x65_c, x71, x78, x81, x82_c, x84, x88_c, x94_c, x96_c, x97, x98_c);
and (w3038, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3039, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3040, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3041, x2_c, x11, x29_c, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3042, x49, x56_c, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3043, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x30, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3044, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x82_c, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3045, x0, x4, x5, x9, x10, x12, x17, x18_c, x19, x20, x22, x25, x26_c, x28, x29_c, x30, x32, x33_c, x34_c, x35_c, x37, x38, x39_c, x40_c, x42, x43_c, x44, x45, x47, x49, x50_c, x51, x52_c, x54, x57_c, x58_c, x59, x61_c, x62_c, x63, x65, x66, x67_c, x68_c, x69, x70, x71, x72_c, x73_c, x74_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85_c, x87, x88_c, x89_c, x91, x92, x93_c, x95, x97, x98_c, x99);
and (w3046, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3047, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3048, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14_c, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3049, x0, x3_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3050, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x46_c, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3051, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75);
and (w3052, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3053, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91_c, x92, x93, x94_c, x95, x96, x98);
and (w3054, x2_c, x11, x29_c, x98_c, x99);
and (w3055, x0, x3, x4, x5, x8_c, x10_c, x12, x13, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3056, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x92_c, x95, x97_c);
and (w3057, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3058, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32_c, x40, x82, x90_c, x96, x98, x99_c);
and (w3059, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3060, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x38, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3061, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3062, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3063, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44, x82, x90_c, x96, x98, x99_c);
and (w3064, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3065, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x58, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3066, x3, x9_c, x14, x34_c, x37, x38_c, x47_c, x60, x67_c, x71, x75_c, x79_c, x81, x82_c, x91, x99_c);
and (w3067, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x39_c, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3068, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x71_c, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3069, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3070, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x77, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3071, x7, x8, x15, x18, x20, x21_c, x26_c, x27, x28, x34, x42, x45_c, x47, x50, x51_c, x52_c, x56_c, x58_c, x69, x71, x76_c, x79, x82, x83_c, x87_c, x92, x94, x96_c, x97_c);
and (w3072, x4, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3073, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x66_c, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3074, x12_c, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3075, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3076, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x47_c, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3077, x2_c, x3_c, x6, x8_c, x11_c, x13_c, x16, x18, x19_c, x24, x25, x26_c, x29_c, x33_c, x34, x35_c, x36, x38_c, x39_c, x40, x44, x45_c, x51, x52_c, x59, x61_c, x67, x76, x80_c, x81, x82_c, x84_c, x85, x86_c, x88, x89_c, x96, x97_c, x98_c);
and (w3078, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3079, x0, x4_c, x15_c, x22_c, x24_c, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3080, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3081, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3082, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x72, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3083, x12_c, x30, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3084, x12_c, x32, x41_c, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3085, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3086, x5_c, x9, x27, x61_c, x76, x78_c, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3087, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3088, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3089, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x51_c, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3090, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x93_c, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3091, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x29_c, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3092, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3093, x0, x1, x2, x4, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3094, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3095, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94, x97_c);
and (w3096, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89_c, x93_c, x95_c);
and (w3097, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x37, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3098, x0, x1_c, x2_c, x3, x4_c, x10, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3099, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x63, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3100, x0_c, x1_c, x2, x3, x5, x6_c, x7, x9_c, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x20_c, x21, x22, x24, x27_c, x29_c, x33, x34_c, x35_c, x36_c, x37, x40_c, x41, x42, x44_c, x45, x46, x49_c, x50, x51_c, x52, x54, x56, x57_c, x58_c, x59, x60, x62_c, x64_c, x65, x69, x70, x71_c, x72_c, x73, x75_c, x77, x78_c, x79, x81, x82, x83, x86_c, x87_c, x89, x91, x92_c, x96_c, x97);
and (w3101, x2, x3, x6_c, x10_c, x11, x13_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3102, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3103, x49, x55_c, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3104, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3105, x0, x4_c, x5_c, x6_c, x7_c, x8_c, x11, x16_c, x18_c, x19, x22, x23, x26, x27, x28, x29, x33, x34, x36, x37_c, x40_c, x41_c, x42_c, x44_c, x46, x47, x49_c, x50, x51, x52_c, x53_c, x54, x56, x57, x60, x61, x63_c, x64, x65_c, x67, x68, x69_c, x70, x72, x75, x76, x77, x79_c, x80_c, x81_c, x83_c, x85, x86_c, x88_c, x91_c, x92, x93, x96, x97, x98_c);
and (w3106, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x98, x99);
and (w3107, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3108, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20_c, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3109, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x87, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3110, x2_c, x3, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3111, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x20, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3112, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x62_c, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3113, x0, x4_c, x15_c, x22_c, x23_c, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3114, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3115, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99_c);
and (w3116, x5, x10, x16, x21_c, x24, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w3117, x0, x2, x3, x6_c, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3118, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x64_c, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w3119, x0, x1, x2_c, x3, x4, x5_c, x6, x7, x8_c, x11_c, x16_c, x17, x18, x19, x20_c, x21, x22_c, x24, x25, x28, x30_c, x31_c, x32_c, x33, x34, x35_c, x36_c, x40_c, x41, x42_c, x43, x44, x45, x46, x47, x48, x50, x51, x52_c, x54, x56_c, x60, x61_c, x63_c, x65_c, x66, x67_c, x68_c, x70, x72, x73, x76, x82, x83_c, x85_c, x86, x88, x89, x92_c, x93_c, x94, x95, x96, x97, x99);
and (w3120, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3121, x0, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3122, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w3123, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x45_c, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3124, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3125, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37, x40, x82, x90_c, x96, x98, x99_c);
and (w3126, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3127, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3128, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3129, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3130, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
assign w3131 = x87_c;
and (w3132, x3_c, x4, x5, x8, x10, x13, x15_c, x17_c, x18, x19_c, x20_c, x21, x23, x24, x25, x27, x30_c, x31, x37_c, x42_c, x44_c, x45_c, x47_c, x49_c, x50_c, x54_c, x55, x58_c, x60, x61_c, x64, x66, x69, x70, x73, x75, x76, x77, x80_c, x81, x83, x86_c, x91, x92, x96, x98, x99);
and (w3133, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3134, x1, x27_c, x35, x36_c, x45, x48, x50, x58, x86_c, x87_c, x92_c);
and (w3135, x4_c, x5_c, x7, x83_c);
and (w3136, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3137, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x26, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3138, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x75_c, x77, x82, x83, x93_c, x95);
and (w3139, x12_c, x32, x69_c, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3140, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x65, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3141, x0_c, x1, x2, x3_c, x4_c, x5, x6, x7, x8, x9, x10, x11_c, x12, x13, x15, x16, x17_c, x18_c, x19, x20_c, x22, x24, x25_c, x26_c, x27_c, x28, x29_c, x30, x31, x32_c, x33, x34, x35, x36_c, x37, x38_c, x40_c, x41, x42, x43, x44_c, x45_c, x46, x47_c, x48, x49, x50_c, x51, x52_c, x53_c, x54_c, x55_c, x57, x59_c, x60, x61_c, x62, x63, x64, x65_c, x66, x67_c, x68_c, x69, x70_c, x71_c, x72, x73_c, x74_c, x75_c, x77, x78, x79_c, x81, x82, x83_c, x84_c, x85_c, x86, x88, x89_c, x90, x91_c, x92_c, x93, x94_c, x96, x97_c, x98, x99);
and (w3142, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3143, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3144, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x69, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3145, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x12_c, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3146, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x75, x84_c, x85_c, x97_c);
and (w3147, x6, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3148, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3149, x5_c, x9, x27, x61_c, x76, x88_c, x92_c, x95, x97_c);
and (w3150, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89, x91);
and (w3151, x0_c, x1, x3, x5_c, x7, x8_c, x9_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3152, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3153, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3154, x4, x5_c, x9_c, x14_c, x15, x18, x19, x20, x21_c, x23_c, x25, x27_c, x30_c, x32, x33_c, x36, x38, x41_c, x46, x47, x48, x49_c, x50_c, x51, x52_c, x53_c, x59, x61_c, x64, x67_c, x69, x71, x75, x78_c, x81, x83_c, x85_c, x87_c, x89_c, x95);
and (w3155, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3156, x13_c, x14_c, x37_c, x39_c, x40_c, x82, x90_c, x96, x98, x99_c);
and (w3157, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17_c, x83_c);
and (w3158, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3159, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3160, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80, x83_c);
and (w3161, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3162, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3163, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61_c, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3164, x13_c, x14_c, x37, x40, x82, x90_c, x96, x98, x99_c);
and (w3165, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3166, x13_c, x49, x64, x71, x72_c, x79, x93, x97_c);
and (w3167, x0_c, x6_c, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3168, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47, x71_c);
and (w3169, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3170, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3171, x3, x8, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3172, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24_c, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3173, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95, x97_c);
and (w3174, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3175, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x38, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3176, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x83_c);
and (w3177, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x14, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3178, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99_c);
and (w3179, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x97, x98, x99_c);
and (w3180, x29_c, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3181, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w3182, x0_c, x4_c, x5_c, x6_c, x8_c, x11_c, x13_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3183, x3_c, x4_c, x5, x7_c, x8_c, x9_c, x11, x14, x15_c, x17_c, x18_c, x21_c, x24, x32_c, x33, x35_c, x40_c, x41, x43_c, x44, x49, x52_c, x53, x59_c, x62, x63_c, x65, x66_c, x70_c, x72_c, x73, x78, x79_c, x82_c, x86, x89_c, x92_c, x93_c, x96, x97, x99);
and (w3184, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x11, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3185, x1, x7, x9, x10_c, x11, x13_c, x14, x15, x17_c, x19, x20_c, x22, x25, x27_c, x29_c, x31_c, x32, x33, x34_c, x39, x40, x43_c, x45, x48, x52_c, x60_c, x61, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x76_c, x78, x79, x82, x83, x84_c, x85, x89_c, x97, x98);
and (w3186, x0_c, x2, x5, x6_c, x9, x11, x12_c, x14, x15, x18, x22, x25, x27_c, x32_c, x35_c, x36, x37, x39, x42, x45_c, x46, x47, x48_c, x50_c, x52, x53, x60_c, x64_c, x67, x68, x70, x71, x75_c, x76, x77_c, x79, x84_c, x87, x91, x98, x99);
and (w3187, x0, x2, x8, x9_c, x10, x13_c, x15_c, x18, x19, x20_c, x21, x23, x24, x25_c, x27, x32, x34, x35, x36_c, x39, x45_c, x49_c, x50, x52, x53_c, x55, x62_c, x64_c, x65, x67_c, x68, x70, x73, x74_c, x75_c, x79_c, x81, x82_c, x83_c, x85_c, x86_c, x88, x92_c, x94_c, x96, x98);
and (w3188, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91, x92_c, x94, x96, x97);
and (w3189, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56_c, x82, x90_c, x96, x98, x99_c);
and (w3190, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3191, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3192, x4_c, x7, x14, x16, x20_c, x25, x31, x32, x42_c, x50, x57_c, x65_c, x71, x74, x75_c, x80_c, x90);
and (w3193, x5, x10, x16, x21_c, x34, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3194, x13_c, x14_c, x20, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3195, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w3196, x1_c, x2, x4, x5_c, x6_c, x8_c, x9, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3197, x1_c, x2, x6_c, x8_c, x14, x17, x21, x22, x28, x32, x33_c, x36, x41, x43_c, x44_c, x46_c, x49, x63_c, x65, x72, x73, x75, x76_c, x87_c, x91_c, x97_c, x99_c);
and (w3198, x0_c, x3_c, x4_c, x6, x7, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3199, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x62_c, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3200, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w3201, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x89_c, x91_c, x92_c, x93, x97_c);
and (w3202, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3203, x4, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3204, x2_c, x5_c, x6, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3205, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94, x95_c);
and (w3206, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3207, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3208, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x90_c, x93_c, x97_c);
and (w3209, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x93_c, x96, x98_c);
and (w3210, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x54, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3211, x0, x2, x3_c, x5, x6_c, x9_c, x12, x13, x14_c, x16_c, x18, x21_c, x24_c, x25, x31_c, x35_c, x37, x40, x41_c, x43, x44_c, x45_c, x46, x47_c, x48, x49_c, x51_c, x52, x54, x55_c, x57_c, x58, x59, x60_c, x63_c, x64, x65, x67, x69_c, x72, x73, x75_c, x77, x78, x80, x82, x84, x88_c, x89_c, x92_c, x93_c, x94, x97, x98, x99);
and (w3212, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88, x89, x93, x97_c, x98_c, x99_c);
and (w3213, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3214, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3215, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3216, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3217, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3218, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3219, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3220, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x71, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3221, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89, x90_c, x91, x92, x95, x97_c);
and (w3222, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x92_c, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3223, x0, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3224, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x60, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3225, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3226, x0, x4, x5_c, x6, x7, x9, x11_c, x12_c, x13_c, x15_c, x16, x18_c, x19, x20, x23_c, x25_c, x26_c, x27_c, x28, x30, x31, x33_c, x35, x39_c, x40_c, x42, x44_c, x48, x49, x50, x51, x53, x54, x57_c, x58, x60, x61_c, x65_c, x66_c, x68, x70, x73, x74, x76_c, x79_c, x80, x81_c, x82, x83_c, x85_c, x86, x87, x88_c, x90, x91_c, x92, x95, x97);
and (w3227, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x95_c, x96_c, x97, x98, x99_c);
and (w3228, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w3229, x0_c, x5, x18, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3230, x2, x4_c, x5, x6, x7_c, x8, x11_c, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3231, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78, x82, x83, x93_c, x97_c);
and (w3232, x1, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3233, x2_c, x11, x29_c, x58, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3234, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x91_c, x95, x96, x97, x99_c);
and (w3235, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3236, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x69, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3237, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8_c, x9_c, x10, x12_c, x13_c, x15_c, x16, x18_c, x19, x21, x23_c, x24, x25, x26, x27, x28_c, x30_c, x31_c, x32, x33, x34_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x45_c, x47_c, x48, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x57_c, x58_c, x60_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80, x82, x83_c, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92_c, x93_c, x94_c, x97, x98, x99_c);
and (w3238, x12_c, x32, x53, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3239, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x28, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3240, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3241, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3242, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86, x93_c, x97_c);
and (w3243, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x21_c, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3244, x1_c, x2_c, x7, x13_c, x18_c, x26, x27_c, x38, x40_c, x51_c, x54_c, x55_c, x61, x63_c, x64, x70_c, x71, x74_c, x82_c, x89_c, x91, x93, x94, x97);
and (w3245, x27, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3246, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x60_c, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3247, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56_c, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3248, x0_c, x2_c, x3_c, x4_c, x6, x7_c, x8, x9_c, x10_c, x11, x12, x13_c, x14, x16, x17, x19_c, x20, x21, x22, x23, x25_c, x27, x31_c, x33, x34, x36_c, x37, x39, x40, x42_c, x43, x44, x45_c, x46_c, x47_c, x48, x49, x50_c, x51_c, x52_c, x55, x56_c, x57, x64_c, x65_c, x66, x67_c, x68, x74, x76, x77_c, x78_c, x79, x80, x81, x84_c, x85, x88_c, x89_c, x93_c, x94_c, x96, x97, x99_c);
and (w3249, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x56_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3250, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98);
and (w3251, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3252, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x93_c, x97_c, x98_c, x99_c);
and (w3253, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3254, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x23, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3255, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x40, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3256, x11_c, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3257, x7, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3258, x0_c, x1, x2, x3_c, x4_c, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x15_c, x17, x18, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26, x27, x28, x29_c, x30_c, x31, x32_c, x33, x34, x35, x36, x37_c, x38_c, x39_c, x40, x41, x42, x43, x45_c, x46, x47, x48, x49, x50, x51, x52, x53, x54_c, x55_c, x56, x57, x59_c, x60_c, x61, x62, x63, x64_c, x65, x66, x67_c, x69_c, x70_c, x71, x72_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80, x81_c, x82, x84_c, x85_c, x86, x87_c, x88_c, x89, x90, x91_c, x92_c, x93_c, x94, x95, x96_c, x97, x98_c, x99_c);
and (w3259, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92_c, x93, x97_c, x98_c, x99_c);
and (w3260, x5, x10, x11, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3261, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3262, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3263, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c, x98_c, x99_c);
and (w3264, x0_c, x1, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3265, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3266, x6_c, x7, x8_c, x11_c, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3267, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x32_c, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3268, x2, x4_c, x5, x6, x7, x8_c, x11_c, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3269, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x12, x40, x82, x90_c, x96, x98, x99_c);
and (w3270, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x62_c, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3271, x2, x6, x8, x11_c, x12_c, x13, x18, x26, x36_c, x42, x43_c, x50, x52_c, x57_c, x61_c, x67, x70, x72_c, x78, x80_c, x82, x86, x88_c, x89_c, x90_c, x95, x97, x99_c);
and (w3272, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x65_c, x66_c, x75_c, x77, x88_c, x93_c, x95_c);
and (w3273, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x30, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3274, x0_c, x3_c, x4_c, x6, x7, x12_c, x40, x82, x90_c, x96, x98, x99_c);
and (w3275, x0_c, x1, x3_c, x4_c, x5_c, x6_c, x7, x8, x9_c, x10_c, x11_c, x12_c, x14, x15_c, x16_c, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25, x26_c, x27_c, x28, x29, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50, x51, x52_c, x54_c, x55_c, x56_c, x57_c, x58_c, x59_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x70, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w3276, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x46, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3277, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x14, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3278, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3279, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3280, x48_c, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3281, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3282, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x63, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3283, x2_c, x3_c, x6, x10, x11, x19, x20_c, x22, x24, x25, x26, x28, x31_c, x33, x34_c, x37, x38_c, x39, x43_c, x45, x46, x50_c, x61, x67, x70_c, x73, x74_c, x76, x81_c, x85, x89, x92_c, x95, x97, x98_c);
and (w3284, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3285, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3286, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x95, x97_c);
and (w3287, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x61, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3288, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3289, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x36_c, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3290, x8, x18_c, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3291, x0_c, x1_c, x3, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3292, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3293, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3294, x8, x9_c, x11_c, x13, x16_c, x17, x18_c, x19, x23, x24, x25, x28_c, x30, x31_c, x33_c, x38, x39, x42, x43, x44, x45, x50, x51_c, x54, x56_c, x59, x63, x68, x69, x72_c, x74_c, x76_c, x79_c, x80_c, x81_c, x84_c, x86_c, x87, x89, x92, x94, x95, x97, x98);
and (w3295, x4_c, x5_c, x7_c, x8_c, x83_c);
and (w3296, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x18, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3297, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3298, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3299, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67, x82, x90_c, x96, x98, x99_c);
and (w3300, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3301, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32_c, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w3302, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3303, x5, x7, x10_c, x11, x12, x15_c, x20_c, x22_c, x27_c, x29_c, x31_c, x35_c, x39, x50_c, x60, x68_c, x71_c, x79, x84_c, x88, x90, x93);
and (w3304, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3305, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x70, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3306, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x36_c, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3307, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x87, x88, x91, x93_c, x97, x98);
and (w3308, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x93_c, x95_c, x96, x98, x99);
and (w3309, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x96, x97, x98, x99_c);
and (w3310, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3311, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3312, x4_c, x33, x44);
and (w3313, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3314, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3315, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x53_c, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3316, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x49, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3317, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3318, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3319, x12_c, x32, x54_c, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3320, x4, x5_c, x6_c, x7, x13, x18_c, x19, x20_c, x21_c, x22_c, x29_c, x33, x34, x35_c, x37, x38, x39_c, x42, x49, x50_c, x51_c, x52, x54, x58_c, x59, x60_c, x63, x66, x67, x70, x71_c, x73_c, x74, x75, x76, x77, x81, x83, x84, x85, x86_c, x93_c, x94_c, x96, x97);
and (w3321, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3322, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3323, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x57_c, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3324, x6, x7_c, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3325, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x75, x77, x82, x83, x93_c, x97_c);
and (w3326, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x66_c, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3327, x0_c, x1_c, x3_c, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3328, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x71_c, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3329, x2_c, x11, x17, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3330, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x38, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3331, x0, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x11_c, x12, x14_c, x15, x17_c, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25, x26, x27, x28_c, x29, x30_c, x31, x32, x33_c, x34_c, x35_c, x36, x37, x38, x40, x41_c, x42, x43_c, x44, x45, x46, x47, x48, x49_c, x50_c, x51, x52, x53_c, x54, x55_c, x56_c, x57_c, x60, x61, x62_c, x63, x65, x66_c, x68, x69_c, x70_c, x71, x72, x73_c, x74, x76_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x85, x86_c, x88, x89, x90, x91, x92, x93, x94, x95, x96_c, x97_c, x98_c);
and (w3332, x11, x12_c, x15, x17_c, x21, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3333, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3334, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x86, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3335, x0_c, x1_c, x2, x3, x4, x6, x7_c, x8, x9_c, x10, x11, x12_c, x13_c, x14_c, x15, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x34, x35, x36, x37, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45_c, x46, x48_c, x49, x50_c, x51_c, x52_c, x53, x54, x56, x57_c, x58_c, x59, x60, x61_c, x62_c, x63_c, x65, x66, x68, x69, x70_c, x71, x72_c, x73, x75, x76, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x86, x87_c, x88, x89, x90, x91, x93_c, x94_c, x95, x96_c, x99_c);
and (w3336, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x73, x76, x85, x89, x93, x97_c);
and (w3337, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x90_c, x93_c, x99_c);
and (w3338, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x89, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3339, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89, x90, x93_c, x97_c);
and (w3340, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3341, x11, x12_c, x15, x17_c, x23_c, x27_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3342, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x83_c, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3343, x6, x7, x11_c, x13, x15_c, x16_c, x17, x18_c, x26_c, x29, x31_c, x33_c, x34_c, x40_c, x41, x43_c, x44, x45, x47, x49_c, x50_c, x51, x52, x58, x59, x64_c, x66_c, x67, x71, x72_c, x75_c, x78, x81_c, x83, x87, x90_c, x91, x92, x94, x95, x96, x98_c, x99_c);
and (w3344, x0_c, x3_c, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3345, x12_c, x32, x91, x97, x98, x99);
and (w3346, x0_c, x1_c, x3, x4_c, x9, x11, x13_c, x20, x23, x24_c, x26_c, x29_c, x30_c, x34_c, x38, x45_c, x46_c, x47_c, x48_c, x49, x51, x52, x56_c, x57, x59_c, x62, x64_c, x69_c, x70_c, x73, x74, x77, x80, x84_c, x89_c, x90, x97, x98_c);
and (w3347, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99);
and (w3348, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x32_c, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3349, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41_c, x83_c);
and (w3350, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x18, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3351, x0, x2, x5_c, x6, x7_c, x8, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3352, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3353, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3354, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3355, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x65, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3356, x0, x2, x3, x6_c, x10_c, x11, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3357, x4_c, x8, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w3358, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x65_c, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3359, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3360, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3361, x12_c, x37_c, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3362, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3363, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x20_c, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3364, x1_c, x4_c, x5, x16, x22_c, x28, x29_c, x33, x38, x41, x42_c, x49_c, x56, x67, x75_c, x81_c, x84_c, x88_c, x91, x94_c, x98_c);
and (w3365, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3366, x0_c, x1, x3_c, x4, x5, x6_c, x7, x8_c, x9_c, x10, x12, x13, x14_c, x16_c, x17, x18_c, x19_c, x20_c, x21, x24, x26, x27_c, x28, x29_c, x32, x35, x36, x37, x45_c, x46, x49_c, x50_c, x52_c, x53, x55, x60, x65_c, x66_c, x67, x68_c, x69, x70_c, x72, x73_c, x75, x76, x78_c, x79_c, x81, x82_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92, x93, x94_c, x97_c, x98, x99);
and (w3367, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3368, x21_c, x26_c, x29, x32_c, x56_c, x79_c, x89_c, x94, x95_c, x97, x98_c);
and (w3369, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3370, x13_c, x49, x64, x71, x72_c, x73_c, x75, x81_c, x87, x90, x93_c, x97_c);
and (w3371, x0, x1, x2, x3_c, x5_c, x6_c, x7_c, x8, x9_c, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x20, x22_c, x23, x24_c, x25_c, x26_c, x27_c, x28, x29, x30_c, x31_c, x33, x34_c, x36_c, x37, x38_c, x39_c, x40_c, x41_c, x42_c, x43, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52_c, x53, x54, x57_c, x58, x59, x60, x61_c, x62, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x76, x77_c, x78_c, x79_c, x80, x81_c, x82, x83_c, x84, x86, x87, x88, x89, x90_c, x91, x92_c, x93, x94_c, x96_c, x97, x98_c, x99_c);
and (w3372, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3373, x1_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3374, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3375, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x57_c, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3376, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74_c, x77, x82, x90_c, x96, x98, x99_c);
and (w3377, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x83_c, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3378, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x48_c, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3379, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3380, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3381, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3382, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3383, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3384, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91, x93_c, x97_c);
and (w3385, x0, x1_c, x5, x6_c, x7, x8, x12, x13_c, x18, x25_c, x33_c, x36, x37_c, x39, x41, x46_c, x48, x49_c, x51_c, x55_c, x62, x68_c, x70, x71_c, x72_c, x74_c, x75, x76, x77, x79_c, x81_c, x86_c, x88_c, x89, x90, x91, x92, x94, x95_c, x98_c);
and (w3386, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3387, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x84_c, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3388, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56, x83_c);
and (w3389, x12_c, x40, x75_c, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3390, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3391, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3392, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9_c, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3393, x23_c, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3394, x69_c, x80_c, x87);
and (w3395, x0, x3, x4, x5, x8_c, x10_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3396, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3397, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3398, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x90_c, x91, x95, x96, x97, x99_c);
and (w3399, x8, x21_c, x25_c, x27_c, x34, x39_c, x44, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3400, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3401, x12_c, x32, x57_c, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3402, x0, x1_c, x2_c, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10, x11_c, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24, x26_c, x27, x28_c, x29, x30, x31, x32_c, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54_c, x56_c, x57, x58_c, x59, x60_c, x61, x62, x63, x64, x65, x66_c, x67, x68_c, x69, x70, x71_c, x72_c, x73_c, x74_c, x75_c, x76, x77_c, x78, x79, x80, x81, x82, x83, x84_c, x85_c, x86, x87, x88, x89_c, x90_c, x91, x92_c, x93_c, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3403, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x97);
and (w3404, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x84, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3405, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3406, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x43, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3407, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37_c, x83_c);
and (w3408, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3409, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3410, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x40, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3411, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84);
and (w3412, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x27_c, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3413, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x13_c, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3414, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37_c, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w3415, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3416, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x55_c, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3417, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74_c, x77_c, x80_c, x82_c, x90_c, x96, x98, x99_c);
and (w3418, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3419, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x58, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3420, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3421, x0, x1_c, x2, x3, x5, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3422, x0, x4_c, x15_c, x22_c, x25_c, x31, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3423, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x87, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3424, x12_c, x32, x64_c, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3425, x0_c, x3_c, x4, x8_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3426, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3427, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x37, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3428, x18, x20_c, x34_c, x51, x58, x75_c, x82, x83_c);
and (w3429, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x40_c, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3430, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3431, x11_c, x43, x53_c, x78, x90_c);
and (w3432, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x79, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3433, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x62_c, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3434, x12_c, x40, x66_c, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3435, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3436, x0, x3, x10, x13, x14, x15, x16_c, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3437, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w3438, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19_c, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3439, x0_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x11, x12_c, x13, x14_c, x15_c, x16, x17, x19, x20_c, x21_c, x22_c, x23, x24_c, x25_c, x26, x27, x28, x29_c, x30, x31_c, x32_c, x33_c, x34_c, x35, x36, x37_c, x38, x39_c, x40, x41, x42, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x54_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63, x64_c, x65, x66_c, x67_c, x68_c, x69_c, x70_c, x71, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79, x80, x81, x82, x83_c, x85, x86, x87_c, x88, x89_c, x90, x92_c, x94, x95_c, x96_c, x97, x98, x99_c);
and (w3440, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x68, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3441, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3442, x1_c, x2, x3, x6_c, x7, x8, x9_c, x11, x15, x16, x18, x19_c, x21, x22, x23, x25, x27_c, x30_c, x31_c, x32, x35, x36_c, x37_c, x38_c, x39_c, x41, x42, x44, x45_c, x46_c, x47, x48_c, x50, x51, x52, x53_c, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61_c, x62, x63_c, x65, x66, x67_c, x68, x70, x71, x73_c, x74, x75, x76, x77, x78_c, x79_c, x81_c, x82_c, x84_c, x87, x88, x92_c, x93_c, x95_c, x96, x97, x98, x99);
and (w3443, x0_c, x3_c, x4_c, x6, x7_c, x11, x13_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3444, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3445, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x74_c, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3446, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3447, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3448, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x55, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3449, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3450, x28_c, x30, x87, x99_c);
and (w3451, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3452, x8, x21_c, x25_c, x27_c, x34, x39_c, x44, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3453, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x95_c, x96, x97_c);
and (w3454, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91_c, x97_c);
and (w3455, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x51, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3456, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3457, x3_c, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3458, x3, x13, x17, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3459, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3460, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3461, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86_c, x93_c, x97_c);
and (w3462, x49, x72, x73_c, x74, x75_c, x79, x90_c, x93_c, x97_c);
and (w3463, x0_c, x5, x23_c, x27_c, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3464, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x49, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3465, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x82_c, x83, x93_c, x97_c);
and (w3466, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x31, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3467, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w3468, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68_c, x73_c, x76, x85, x89, x93, x97_c);
and (w3469, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3470, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89, x90_c, x91_c, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3471, x0, x1, x2, x3_c, x4, x5, x6, x7, x8, x9, x10_c, x11, x12_c, x13, x14_c, x15_c, x16, x17, x18_c, x19_c, x20, x21_c, x22_c, x23, x25_c, x26_c, x27_c, x28_c, x29, x30_c, x31, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x40_c, x41_c, x43, x44, x45_c, x48_c, x50_c, x51_c, x52, x53, x54, x55_c, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x67_c, x68, x69_c, x70_c, x71, x72_c, x73, x74_c, x76_c, x77_c, x78_c, x79, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x89, x90_c, x91, x93_c, x94_c, x95, x96_c, x97, x98_c, x99);
and (w3472, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3473, x49, x77_c, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3474, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3475, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3476, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x19_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3477, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3478, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x45_c, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3479, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x35_c, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3480, x5, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3481, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3482, x49, x69_c, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3483, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x88, x90_c, x91, x92, x95, x97_c);
and (w3484, x11_c, x15_c, x16, x18, x21_c, x23_c, x71_c);
and (w3485, x1_c, x3_c, x6, x9, x10, x13, x14_c, x17_c, x18, x19, x21_c, x22_c, x23_c, x24_c, x27, x28_c, x29_c, x30, x31_c, x36, x38_c, x39_c, x40_c, x41, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x52, x54, x57_c, x58, x59, x60, x62, x64_c, x67, x68_c, x70_c, x72, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81_c, x82, x84_c, x87_c, x89, x90, x92_c, x93, x94_c, x96_c, x97, x98);
and (w3486, x1_c, x2_c, x3, x4, x5, x7, x9, x10_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3487, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98_c);
and (w3488, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3489, x19, x26_c, x34, x35, x38_c, x40, x44, x59, x60, x68, x78, x86_c, x87_c, x99_c);
and (w3490, x1_c, x4, x8, x33_c, x44_c, x69, x81, x85, x91, x97_c);
and (w3491, x0_c, x5, x10_c, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3492, x1_c, x2_c, x6, x8, x9_c, x10_c, x12_c, x14, x16_c, x17, x18_c, x19, x20, x21_c, x22_c, x24_c, x25, x26, x30, x31_c, x34, x35_c, x36_c, x37_c, x39, x41_c, x45_c, x46_c, x50, x51, x52_c, x61, x63, x64_c, x66, x68, x69_c, x71, x72, x75, x76_c, x78, x79, x80_c, x82, x84_c, x85, x88_c, x89_c, x94_c, x96, x97, x98_c, x99_c);
and (w3493, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x32, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3494, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x71_c, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3495, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3496, x0, x1_c, x2_c, x4_c, x5, x16, x17, x18, x19, x20_c, x21_c, x22_c, x24_c, x25, x27_c, x28_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x36_c, x38, x40_c, x43, x44, x45, x46, x47, x51_c, x52_c, x53_c, x54, x56_c, x58_c, x61, x62, x64_c, x65, x66, x68_c, x71_c, x72, x73, x74_c, x76_c, x77, x81, x87, x89, x91, x94_c, x95_c, x96, x99);
and (w3497, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x34, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3498, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3499, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25_c, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3500, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3501, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x69, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3502, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92, x93, x94_c, x96_c, x97_c, x98_c, x99);
and (w3503, x1, x3, x4, x6_c, x8_c, x11_c, x14, x15, x20_c, x22_c, x23, x24, x25, x26, x27_c, x30_c, x31_c, x33, x34_c, x35, x36_c, x37, x38, x39, x41_c, x43, x44_c, x48, x49_c, x50, x51, x53_c, x55_c, x56_c, x58, x59, x60_c, x62, x63, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x73_c, x74, x76, x78_c, x80_c, x82_c, x83, x84, x85, x86, x87_c, x89_c, x90_c, x91_c, x93_c, x96, x97_c);
and (w3504, x3, x9_c, x11_c, x19, x24_c, x27_c, x35_c, x39, x55, x56_c, x72, x89_c);
and (w3505, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54, x73_c, x76, x85, x89, x93, x97_c);
and (w3506, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72_c, x83_c);
and (w3507, x8, x21_c, x25_c, x27_c, x34, x38, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3508, x0, x3_c, x5, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3509, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x86_c, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3510, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x47_c, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w3511, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43_c, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3512, x3_c, x4, x5, x6, x7_c, x9, x12_c, x13, x14, x15, x18, x24_c, x27_c, x31, x32, x34, x36_c, x38, x40_c, x44, x48_c, x49, x53, x56_c, x57, x58, x59, x60, x61, x62, x65, x66_c, x67, x70, x71_c, x73_c, x75_c, x76_c, x78, x81, x83, x85, x87_c, x88_c, x94, x95, x96_c);
and (w3513, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3514, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3515, x12_c, x32, x34_c, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3516, x49, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3517, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73_c, x83_c);
and (w3518, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3519, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3520, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3521, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3522, x6, x17_c, x20_c, x24_c, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w3523, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x82, x90_c, x96, x98, x99_c);
and (w3524, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3525, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x36_c, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3526, x0_c, x1, x2, x5_c, x6, x7_c, x10, x13_c, x14, x16, x17_c, x22, x24_c, x26, x29, x30_c, x32, x35, x37, x38_c, x39_c, x40_c, x43_c, x44_c, x45_c, x47, x48_c, x50, x54_c, x56_c, x58_c, x59, x60_c, x61_c, x62, x65, x67, x68, x71, x73_c, x76_c, x80_c, x81, x83_c, x84, x85_c, x88, x89_c, x90_c, x92_c, x96);
and (w3527, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3528, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3529, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3530, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3531, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3532, x5_c, x9, x27, x60, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3533, x5, x10, x16, x21_c, x28, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w3534, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x61, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3535, x3_c, x5, x6_c, x9, x10_c, x14_c, x15_c, x24, x25, x27, x29_c, x31, x32_c, x34, x35_c, x37, x38, x41, x43, x44_c, x46, x48, x50, x51, x53_c, x54, x57_c, x58_c, x62, x63_c, x68_c, x69_c, x71_c, x72, x73, x77, x78_c, x79_c, x80, x82_c, x83_c, x84_c, x85, x86_c, x88_c, x90_c, x92, x93);
and (w3536, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x29, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3537, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3538, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x16_c, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3539, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3540, x0, x1_c, x2_c, x3, x4_c, x5_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23, x24, x25_c, x26, x27, x28, x29, x30, x31, x32_c, x33_c, x34_c, x35, x36_c, x37, x38_c, x39_c, x40, x41_c, x42, x43_c, x44_c, x45, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57_c, x58, x59, x60, x61_c, x62, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78, x79, x80, x81, x82_c, x83_c, x84, x85_c, x86, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x97, x98, x99);
and (w3541, x12_c, x20, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3542, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3543, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3544, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x74_c, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3545, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x74_c, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3546, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3547, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3548, x2_c, x3, x4, x5_c, x6_c, x7, x9, x12, x13_c, x14, x15, x16, x17, x18, x19_c, x21, x23_c, x25_c, x26_c, x27, x28, x29, x30_c, x32, x33, x34, x35, x36_c, x37_c, x38, x39, x40, x41, x42, x43_c, x44_c, x45, x46_c, x47, x48_c, x49, x50_c, x51_c, x52_c, x53_c, x54, x56, x57_c, x59_c, x60, x61, x62_c, x63_c, x64_c, x65, x66_c, x68_c, x69, x70, x71, x72, x74_c, x75, x76, x77, x78_c, x79, x80, x81_c, x83, x85, x86_c, x87_c, x88, x89_c, x90, x91, x94, x96_c, x97, x98_c, x99);
and (w3549, x41_c, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3550, x0, x1, x2, x4, x8_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3551, x0, x3, x10, x13_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3552, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x19, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3553, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3554, x22, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3555, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3556, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x33, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w3557, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x35, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3558, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3559, x10_c, x35, x49_c, x64_c, x95_c);
and (w3560, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x96, x97_c, x98, x99_c);
and (w3561, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3562, x0, x1, x2, x4_c, x5_c, x6_c, x7, x11_c, x12_c, x13, x15, x16_c, x17_c, x18, x19, x20, x23_c, x24, x26, x28_c, x29_c, x30_c, x31, x32, x34_c, x35_c, x36_c, x37, x38, x39_c, x41, x42_c, x43, x46_c, x47_c, x48, x50_c, x51_c, x52, x53_c, x54, x56, x57_c, x58_c, x60, x61_c, x63, x64_c, x65, x66, x67, x68_c, x71_c, x72, x74, x75_c, x76_c, x77_c, x79_c, x83, x84_c, x86_c, x87, x88, x89, x91_c, x92_c, x94, x95, x96_c, x98, x99_c);
and (w3563, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3564, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30_c, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3565, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3566, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3567, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3568, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3569, x0_c, x1_c, x2_c, x4, x6, x7, x8_c, x9, x11_c, x13_c, x17, x18, x19, x20, x22, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x35_c, x36, x38, x39, x41_c, x42_c, x43_c, x44, x45, x46_c, x47_c, x48_c, x49, x50_c, x53, x54, x55, x56_c, x57_c, x58, x60_c, x62, x65_c, x67, x68, x69, x72, x74_c, x76_c, x78, x79, x81, x82_c, x84, x85, x86_c, x87_c, x88_c, x90_c, x91, x92, x94, x95_c, x96_c, x99);
and (w3570, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x70_c, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3571, x0, x3, x10, x13, x14, x15, x16_c, x22, x29_c, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3572, x9_c, x10_c, x12, x15_c, x16, x25_c, x26_c, x27_c, x34, x36, x37, x39_c, x42_c, x56_c, x59_c, x86_c, x88, x93, x95, x98_c);
and (w3573, x1, x2_c, x6, x7_c, x8, x9, x10_c, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3574, x0, x2_c, x4_c, x15_c, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3575, x12_c, x21_c, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3576, x25, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3577, x0, x1, x2_c, x3, x4, x6_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3578, x0_c, x2, x5, x8, x12_c, x14_c, x18_c, x22_c, x24_c, x25_c, x27, x33, x40_c, x47_c, x48, x52, x54_c, x55_c, x61, x62, x63, x70_c, x74_c, x79_c, x80, x84, x85_c, x86_c, x87, x89_c, x91, x92_c, x93_c, x94, x95_c, x96, x99);
and (w3579, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3580, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3581, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3582, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3583, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91_c, x93_c, x97_c);
and (w3584, x5_c, x8, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3585, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x75_c, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3586, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3587, x6_c, x17, x25_c, x38, x48_c, x58_c, x66_c, x68_c);
and (w3588, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3589, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x35_c, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3590, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3591, x0_c, x2_c, x4, x5, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3592, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x19, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3593, x12_c, x40, x64_c, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3594, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x55_c, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3595, x2, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3596, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3597, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3598, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3599, x0_c, x1_c, x2, x4, x5, x6, x7_c, x9_c, x10_c, x11, x12, x13, x14_c, x15_c, x16, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24, x25_c, x27_c, x28, x29_c, x30, x32_c, x33, x37_c, x39, x40_c, x41_c, x43_c, x45_c, x47_c, x48_c, x49, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59, x60, x61, x62_c, x63, x64_c, x65_c, x66_c, x68_c, x69_c, x70, x71, x73, x74_c, x77_c, x78_c, x80, x81_c, x82, x83, x84, x85_c, x86, x88, x90_c, x91_c, x95, x96, x97, x98_c);
and (w3600, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3601, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3602, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3603, x13_c, x47_c, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w3604, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3605, x5, x7, x15_c, x23_c, x29_c, x38_c, x39, x40, x42, x44_c, x52, x53, x59_c, x65_c, x66, x74, x77_c, x81, x82, x87_c, x97);
and (w3606, x8, x21_c, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3607, x0_c, x1, x4_c, x5_c, x6_c, x9_c, x13, x18, x19_c, x24_c, x26, x27_c, x28_c, x29_c, x34_c, x35_c, x36_c, x38, x39, x42, x43_c, x44, x45, x46, x47, x49_c, x54, x56_c, x58, x59_c, x60, x61_c, x63, x64_c, x65_c, x66_c, x71, x73_c, x74_c, x75, x77_c, x78_c, x79, x81_c, x82, x84_c, x86_c, x87, x88_c, x89_c, x91, x93_c, x94_c, x95_c, x96_c, x98);
and (w3608, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x24, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3609, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3610, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x78, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3611, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3612, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x63, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3613, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3614, x5, x10, x16, x17, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w3615, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3616, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3617, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x42, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3618, x0, x1_c, x2_c, x3, x4, x5, x6, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3619, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92, x95);
and (w3620, x10, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3621, x2_c, x11, x29_c, x45, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3622, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x57_c, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3623, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x91_c, x92, x95, x97_c);
and (w3624, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3625, x0, x1, x2_c, x3, x4, x6, x7, x8_c, x9_c, x11_c, x12, x13, x14, x15_c, x17, x18, x19_c, x20, x21, x22_c, x23, x24, x25, x26, x27, x28, x29_c, x30, x31_c, x33_c, x34, x36_c, x37_c, x39, x40, x41, x42, x43, x44_c, x45_c, x46, x47, x48_c, x49, x50, x51_c, x52_c, x53_c, x54, x55_c, x56, x57, x58, x59_c, x60_c, x61_c, x62, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x80, x81_c, x82_c, x83_c, x84_c, x86_c, x87, x88_c, x89, x90_c, x92, x93_c, x94_c, x96, x97_c, x98, x99);
and (w3626, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3627, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3628, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x50, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3629, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91_c, x93_c, x97_c);
and (w3630, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x23, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3631, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w3632, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x69_c, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3633, x6, x8_c, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3634, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3635, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x23, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3636, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x69_c, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3637, x49, x81_c, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3638, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3639, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x72, x79, x90_c, x93_c, x97_c);
and (w3640, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x34_c, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3641, x0_c, x1, x2_c, x3, x4, x7, x8_c, x9, x10, x11, x12, x13_c, x14_c, x15, x16_c, x17_c, x18, x19_c, x20_c, x21, x22_c, x23, x24_c, x25_c, x26_c, x28, x29, x30_c, x31_c, x32, x33, x34, x35, x36, x37, x38, x39_c, x40, x41_c, x43, x44_c, x45_c, x47_c, x48_c, x49, x50, x51_c, x52_c, x53, x54_c, x55, x56, x57_c, x59, x60_c, x61, x63, x65, x66_c, x67, x69, x70, x71, x72_c, x73, x74, x76_c, x77, x78, x80, x81, x83_c, x84, x85_c, x86, x87, x88, x89_c, x90, x91, x92, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w3642, x12_c, x32, x76, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3643, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87_c, x88, x89_c, x90_c, x91_c, x92, x93, x95, x96_c, x97_c);
and (w3644, x0, x3, x10, x13, x14, x15, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3645, x3, x14, x21, x23_c, x24_c, x32_c, x33, x37_c, x38, x45, x59, x61, x70_c, x76_c, x77, x84_c, x87_c, x89, x92);
and (w3646, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3647, x12_c, x28, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3648, x6, x7, x10, x17, x20_c, x22, x33_c, x45, x46, x50_c, x54, x62, x64, x66_c, x68_c, x71, x73, x74_c, x77, x79, x84, x86_c, x90, x96, x97_c, x99);
and (w3649, x12_c, x13_c, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3650, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43_c, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3651, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x21, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3652, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3653, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x66_c, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3654, x13, x14, x23, x24_c, x29_c, x30_c, x42, x43_c, x45, x53_c, x55_c, x56, x64_c, x76_c, x80);
and (w3655, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49, x83_c);
and (w3656, x0, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3657, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3658, x73, x90, x93_c, x95_c, x96, x98, x99);
and (w3659, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3660, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x78_c, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3661, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x89, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3662, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x78, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3663, x4_c, x14_c);
and (w3664, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x48_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3665, x0, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3666, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39, x83_c);
and (w3667, x8, x21_c, x25_c, x27_c, x29_c, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3668, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3669, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3670, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x68, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3671, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3672, x26, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3673, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3674, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3675, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x91, x92_c, x94_c, x96_c, x97_c, x99_c);
and (w3676, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91, x92, x93_c, x94_c, x96, x98, x99);
and (w3677, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3678, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x81_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3679, x4, x6_c, x7, x8, x9, x10, x18, x25, x28, x31_c, x34, x36, x37_c, x38, x40, x41_c, x42_c, x43_c, x45, x46_c, x56_c, x58_c, x60, x62, x64, x69_c, x71, x72_c, x73_c, x77, x78, x81_c, x83, x85, x89_c, x90_c, x93, x94_c, x96, x99);
and (w3680, x0_c, x1, x2_c, x5, x6_c, x7_c, x9_c, x10, x11, x12_c, x13, x14, x15, x16_c, x17, x19_c, x20, x21_c, x22_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x36_c, x37, x38, x39_c, x40, x41_c, x42, x43_c, x44_c, x45_c, x46, x47, x48_c, x49_c, x50_c, x52_c, x53_c, x54_c, x55, x56, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x76, x77, x78_c, x79_c, x80_c, x81_c, x82, x83, x84_c, x85_c, x86, x87_c, x89, x90, x91, x92_c, x93, x94, x95_c, x96_c, x98_c, x99);
and (w3681, x0, x1_c, x2, x9, x11, x12, x20, x23_c, x27_c, x29, x32, x33, x41, x47, x48_c, x49, x50_c, x51_c, x52, x55, x56, x59_c, x60_c, x61_c, x62, x64_c, x69, x71_c, x73, x74, x77_c, x86_c, x89, x91, x99);
and (w3682, x1_c, x2, x3, x4, x5_c, x8, x9_c, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3683, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x95, x96_c, x97_c, x98, x99_c);
and (w3684, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92_c, x93_c, x97_c);
and (w3685, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3686, x5_c, x7_c, x10, x13, x14_c, x16, x19, x20_c, x21_c, x22, x25, x27, x33, x42_c, x45, x47_c, x48, x49_c, x54_c, x58_c, x60, x66_c, x71, x72_c, x73_c, x77_c, x82_c, x85_c, x86, x87, x91, x92, x94, x95);
and (w3687, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3688, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x53_c, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3689, x0_c, x5_c, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3690, x3, x13_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3691, x5_c, x9, x27, x61_c, x76, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3692, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13_c, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3693, x11, x12_c, x15, x17_c, x23_c, x27, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3694, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x22_c, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3695, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3696, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x35, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3697, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3698, x0, x3_c, x4, x6_c, x7, x8, x9_c, x11_c, x12, x13_c, x15, x17, x18_c, x19_c, x22_c, x23, x24_c, x25_c, x26, x28, x30, x31_c, x33_c, x35, x38, x40, x42_c, x43_c, x45, x46_c, x47, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x55, x57_c, x58, x59, x60, x61_c, x62, x64_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x72, x73_c, x74, x75, x76_c, x77, x80, x81_c, x83_c, x84, x88, x90_c, x92_c, x95_c, x98_c);
and (w3699, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3700, x0_c, x1, x2, x3_c, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3701, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3702, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c, x99);
and (w3703, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x52_c, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3704, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x59_c, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3705, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3706, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x24, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3707, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81, x85, x89, x93, x97_c);
and (w3708, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x34_c, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3709, x73, x93, x95_c, x96, x98, x99);
and (w3710, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3711, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3712, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x51_c, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3713, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3714, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x90_c, x93_c, x94, x95, x96, x97_c, x98, x99);
and (w3715, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3716, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3717, x0, x3, x10, x13, x14, x15, x16_c, x22, x34_c, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3718, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x47, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3719, x0, x1, x2_c, x3_c, x8_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3720, x10_c, x16_c, x19, x29_c, x31, x33_c, x34, x42_c, x48_c, x54_c, x60_c, x64_c, x75_c, x85, x88_c, x89, x98, x99);
and (w3721, x1, x4_c, x6, x8, x11_c, x12_c, x15_c, x17, x20_c, x21_c, x24, x27_c, x28, x37, x39_c, x41_c, x43_c, x47, x49, x50, x52_c, x53_c, x57_c, x62_c, x69_c, x73, x76_c, x81, x82_c, x86, x88_c, x89_c, x90, x91_c, x93, x94, x95);
and (w3722, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76_c, x83_c);
and (w3723, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57_c, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3724, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x78_c, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3725, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3726, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x21, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3727, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x61, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3728, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x16_c, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w3729, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3730, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x31_c, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3731, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3732, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3733, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31_c, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3734, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3735, x2_c, x11, x29_c, x36_c, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3736, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3737, x0, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3738, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x68_c, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3739, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3740, x1, x2, x4, x15_c, x18_c, x19_c, x21, x26_c, x28_c, x29_c, x38, x39_c, x47_c, x48, x49_c, x53_c, x58, x59, x62_c, x77, x79, x80, x82_c, x86_c, x87);
and (w3741, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92, x93_c, x95_c, x96);
and (w3742, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44, x83_c);
and (w3743, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x82, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3744, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3745, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x70_c, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3746, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x67_c, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3747, x1_c, x2, x4, x6_c, x7, x8, x10, x12, x18, x20, x21, x22_c, x23_c, x24, x25_c, x26_c, x27_c, x30, x31_c, x32_c, x36_c, x39, x42_c, x44_c, x46, x47_c, x48, x49_c, x51_c, x54_c, x55, x56, x57, x58_c, x66, x69_c, x71, x72, x75_c, x79, x82_c, x83, x84_c, x85, x88, x89_c, x90_c, x92_c, x95, x96_c);
and (w3748, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x55, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3749, x11, x12, x18, x20, x23_c, x26, x29, x41_c, x63, x65, x70, x71_c);
and (w3750, x5, x10, x16, x21, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3751, x0, x1, x2, x3, x5, x6_c, x7, x8, x9_c, x10_c, x11_c, x12_c, x13_c, x14, x15, x16, x18, x19, x20, x21, x22_c, x23, x24, x26, x27_c, x28_c, x29, x32_c, x33_c, x35_c, x36, x37, x38, x39_c, x41, x43, x44, x45_c, x46, x47_c, x48, x49_c, x52, x54, x56_c, x58, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72_c, x73, x74_c, x75_c, x76_c, x78_c, x79, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x88, x89_c, x90_c, x91, x92, x93_c, x94, x95, x96_c, x97, x99_c);
and (w3752, x0, x37, x49, x85_c);
and (w3753, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96_c, x97_c);
and (w3754, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3755, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3756, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3757, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3758, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3759, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89, x90_c, x93_c, x97_c);
and (w3760, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x69, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3761, x0, x1_c, x2, x3, x4, x5, x6_c, x7, x8_c, x9_c, x10, x11_c, x13_c, x14, x15_c, x16, x17_c, x19_c, x20_c, x22_c, x23, x24_c, x25, x26_c, x28, x29_c, x30, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37, x38, x39_c, x40, x41_c, x43, x44, x45, x46, x47_c, x48, x49_c, x50_c, x51_c, x52, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61, x62, x63, x64, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84, x85_c, x86, x87, x89, x90, x91, x92_c, x93, x94_c, x95, x96, x97_c, x98, x99_c);
and (w3762, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3763, x0, x3, x10, x13, x14, x15_c, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3764, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3765, x12_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3766, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3767, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3768, x0_c, x3_c, x4, x12_c, x40, x82, x90_c, x96, x98, x99_c);
and (w3769, x13, x20_c, x21, x26, x30_c, x31, x36, x39, x40, x43, x44_c, x47, x59_c, x68, x71_c, x76, x80, x81, x86_c, x87, x88_c, x99);
and (w3770, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x93_c, x95_c, x97, x99);
and (w3771, x0, x1, x2_c, x3_c, x5_c, x9_c, x11, x16, x19_c, x21, x25, x26_c, x27, x28, x30, x32, x33, x34_c, x35_c, x36_c, x37_c, x39, x41_c, x44, x45, x46_c, x50, x51_c, x52, x54_c, x55_c, x56_c, x57_c, x58_c, x60_c, x61_c, x63_c, x64, x66, x67_c, x70, x71_c, x75_c, x79_c, x80, x81, x82_c, x84_c, x88_c, x90, x91_c, x92, x94, x96, x98_c);
and (w3772, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3773, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24_c, x83_c);
and (w3774, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x74_c, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3775, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3776, x0, x4_c, x15_c, x17_c, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3777, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3778, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x52, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3779, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x84_c, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3780, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3781, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73_c, x74_c, x77_c, x80, x82, x90_c, x96, x98, x99_c);
and (w3782, x2, x3, x6, x7, x8, x9, x12_c, x14_c, x16, x17, x24_c, x25_c, x26_c, x29, x32, x34_c, x35_c, x39_c, x40_c, x41_c, x42_c, x48_c, x49_c, x50, x53, x55, x56_c, x62, x63_c, x64, x65, x69_c, x70, x71_c, x72, x74, x75_c, x76_c, x77, x80_c, x81_c, x83_c, x84, x85_c, x88, x91, x92, x94_c, x96, x97, x98);
and (w3783, x12_c, x30, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3784, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3785, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x42_c, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3786, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3787, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3788, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65, x71_c);
and (w3789, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3790, x1_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17, x18, x19, x20_c, x21_c, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32, x33, x34_c, x35, x36_c, x37, x38, x39, x40, x41, x42_c, x43, x44, x45, x46, x47, x48, x49_c, x50_c, x51, x52, x53_c, x54, x55_c, x56_c, x57_c, x58_c, x59_c, x60, x61, x62, x63, x64_c, x65, x66, x67, x68_c, x69, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78, x79_c, x80, x82, x83_c, x85_c, x86_c, x87_c, x88, x89, x90, x92_c, x93_c, x94, x95_c, x96, x97, x98);
and (w3791, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80, x82, x83, x93_c, x97_c);
and (w3792, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x54_c, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3793, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x40, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3794, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3795, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x56_c, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3796, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3797, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13_c, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3798, x0, x4, x31, x36, x41, x47_c, x54_c, x77_c, x80, x84_c, x87_c, x95_c, x96_c);
and (w3799, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3800, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3801, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3802, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3803, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52_c, x83_c);
and (w3804, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3805, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81_c, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3806, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91, x92_c, x94, x96_c, x97_c);
and (w3807, x0, x1_c, x2, x3, x4, x6_c, x7_c, x8, x9, x10_c, x11_c, x12, x15_c, x18, x20, x21, x23, x27_c, x28_c, x30_c, x37, x41_c, x42_c, x44, x46_c, x49, x57, x60_c, x61_c, x64, x66, x71_c, x72, x73_c, x76_c, x77_c, x78, x82, x83_c, x95_c, x96, x97_c, x98, x99_c);
and (w3808, x0_c, x1_c, x2_c, x3, x5_c, x6, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3809, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3810, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x65_c, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3811, x4_c, x6_c, x12_c, x14, x20_c, x23, x31, x32, x33, x38, x39_c, x40, x42_c, x43_c, x44, x48, x53, x56, x58_c, x59, x60, x61, x63_c, x64_c, x66, x70, x72, x74, x75, x77, x78, x80_c, x82, x84_c, x87, x88, x94);
and (w3812, x0, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3813, x1_c, x3_c, x4, x6_c, x13_c, x21_c, x23, x24_c, x33, x37, x46, x49_c, x54, x55, x57, x58_c, x59, x61, x63, x68_c, x80, x81_c, x89_c, x91_c, x95);
and (w3814, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x63, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3815, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3816, x3_c, x9_c, x15_c, x18_c, x19_c, x24_c, x26, x28, x29_c, x30, x31, x33_c, x36, x39_c, x41, x42_c, x43, x45, x49, x56_c, x57_c, x58_c, x59_c, x61, x62, x63_c, x71_c, x74, x77_c, x80, x81_c, x82, x83_c, x91_c, x93_c, x94_c, x95, x97, x98_c);
and (w3817, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3818, x13_c, x36, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w3819, x0, x1, x3, x5_c, x7_c, x8_c, x10_c, x11, x12_c, x13, x17, x18_c, x19, x21_c, x22, x23, x25, x30_c, x34_c, x35_c, x36_c, x37_c, x39_c, x42_c, x43, x44_c, x45, x46_c, x49_c, x51_c, x52_c, x53, x57, x59, x60_c, x61_c, x64_c, x68, x69, x70_c, x72_c, x73, x74_c, x75, x76_c, x79, x81, x84_c, x88, x89_c, x92_c, x93_c, x96);
and (w3820, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88, x89_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3821, x1, x2_c, x4_c, x5_c, x7_c, x8, x9, x11_c, x12, x13_c, x16_c, x18, x20_c, x21_c, x22, x23, x24, x27_c, x29, x31, x32_c, x33, x36_c, x37, x38_c, x39, x40, x41, x42, x44, x45, x46, x47_c, x48_c, x49_c, x53_c, x54_c, x55_c, x57_c, x58, x61_c, x63, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71, x72, x73, x75_c, x76_c, x77_c, x78_c, x79, x81_c, x83_c, x84_c, x88_c, x90, x91_c, x92_c, x94_c, x95_c, x98_c, x99);
and (w3822, x39_c, x88_c);
and (w3823, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3824, x9_c, x17_c, x26_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3825, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x92_c, x94_c, x95_c, x96, x97_c);
and (w3826, x5, x6_c, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w3827, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x83_c);
and (w3828, x0, x1, x3, x4_c, x5_c, x7, x8, x9, x12_c, x13, x14_c, x15, x17_c, x18, x19_c, x20, x22, x23, x24_c, x25, x26_c, x28_c, x29, x30, x33, x34, x35, x36_c, x37, x38_c, x39, x40, x42_c, x43, x45_c, x47, x48, x51, x52, x53, x55_c, x56_c, x57, x58, x59_c, x61_c, x65_c, x66_c, x67_c, x68_c, x72, x73_c, x74, x76, x77_c, x78, x81, x82, x83, x84_c, x85, x88, x90, x91_c, x92, x93_c, x95_c, x96_c, x97, x98, x99_c);
and (w3829, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3830, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3831, x49_c, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3832, x8, x21_c, x24, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3833, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3834, x0, x1, x2, x3, x5_c, x8_c, x9_c, x11, x12_c, x13, x14_c, x16, x18_c, x19_c, x20, x21_c, x22, x23, x24, x25_c, x26_c, x27, x28, x29, x30, x31_c, x32_c, x36_c, x37_c, x39_c, x41, x42_c, x43_c, x45, x47, x48, x49, x50, x51_c, x52_c, x54_c, x55, x58, x60_c, x62, x64, x65_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75, x76_c, x77_c, x79, x80_c, x81, x83_c, x84_c, x85, x86, x88, x89_c, x91_c, x92_c, x93_c, x94, x95, x96_c, x97_c);
and (w3835, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3836, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x87_c, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3837, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62_c, x83_c);
and (w3838, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97, x98_c, x99_c);
and (w3839, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3840, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49_c, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3841, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x20, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3842, x3_c, x8, x13_c, x15, x17_c, x27, x28_c, x29, x31_c, x38_c, x40, x42, x43_c, x44_c, x46_c, x49, x52_c, x53, x56_c, x57_c, x58_c, x60, x63_c, x69, x75_c, x76_c, x77_c, x79, x84, x85_c, x92_c, x98);
and (w3843, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x97_c);
and (w3844, x6, x26_c, x34_c, x41, x44_c, x49_c, x60, x71, x77_c, x90_c, x93_c);
and (w3845, x5, x10, x16, x21_c, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3846, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3847, x4_c, x10, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w3848, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x51_c, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w3849, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3850, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3851, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x41_c, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3852, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3853, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x97_c);
and (w3854, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3855, x5_c, x9, x12_c, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3856, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3857, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57_c, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3858, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x55, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3859, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3860, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3861, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3862, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x74, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3863, x0_c, x1, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3864, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57_c, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3865, x0, x1_c, x3, x4_c, x5, x9_c, x12, x16_c, x18, x20_c, x21, x22, x23, x25, x26_c, x27, x28, x32, x36, x37_c, x38, x40, x45, x48_c, x49, x50_c, x51_c, x55, x56, x57_c, x59, x60, x67, x68_c, x69_c, x71, x72_c, x77_c, x78, x80, x81_c, x82_c, x83, x85_c, x87_c, x88, x90, x91_c, x93, x94_c, x98, x99);
and (w3866, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3867, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3868, x49, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3869, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3870, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3871, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48_c, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w3872, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x32_c, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3873, x6, x17_c, x20_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3874, x49, x64, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3875, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3876, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x81_c, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3877, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3878, x3_c, x6, x7, x22_c, x25_c, x28_c, x32, x35, x37, x40, x45_c, x46, x47_c, x50, x56, x63_c, x66_c, x67_c, x69, x71, x75, x81_c, x84, x92_c);
and (w3879, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x36_c, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3880, x0_c, x1_c, x3, x4_c, x5_c, x6, x7, x8, x10_c, x11_c, x12, x13_c, x14, x16_c, x17, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x25, x26_c, x27, x28, x29, x31, x32, x33, x35_c, x37, x38, x40_c, x42_c, x43_c, x44_c, x45_c, x46, x48, x52, x56_c, x58, x59, x60, x61, x62, x63, x64, x65, x66_c, x67_c, x69_c, x70, x71, x72, x73, x74, x75, x76_c, x78_c, x79_c, x81_c, x82, x83, x84, x85_c, x86, x88_c, x89_c, x90_c, x92_c, x93, x96_c, x97_c, x99);
and (w3881, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3882, x1_c, x4_c, x13_c, x14_c, x15, x33, x35, x38_c, x39_c, x40, x41, x46, x48, x50, x51_c, x52, x54, x56, x57_c, x58, x63_c, x64, x68, x70, x71, x72, x76, x78_c, x86_c, x88_c, x96, x99);
and (w3883, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98);
and (w3884, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x62, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3885, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3886, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x86, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3887, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3888, x8, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3889, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3890, x8, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3891, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x41, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3892, x5_c, x9, x27, x58_c, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3893, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3894, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79, x80_c, x82, x83_c, x84_c, x91);
and (w3895, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x95_c);
and (w3896, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3897, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x42, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3898, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3899, x17, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3900, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3901, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3902, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x64_c, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3903, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3904, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3905, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3906, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3907, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13_c, x40, x82, x90_c, x96, x98, x99_c);
and (w3908, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3909, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3910, x0, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3911, x0, x12_c, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3912, x13, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3913, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3914, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x60_c, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3915, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3916, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3917, x0_c, x5_c, x6, x12_c, x13_c, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3918, x0, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3919, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x11, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3920, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91_c, x92, x93, x94_c, x96, x98, x99_c);
and (w3921, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x57, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w3922, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3923, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3924, x0, x1_c, x2, x3, x10, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3925, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3926, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x70, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w3927, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x94_c, x95_c);
and (w3928, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x59_c, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3929, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3930, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92_c, x94_c, x95_c, x97_c);
and (w3931, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78_c, x79, x90_c, x93_c, x97_c);
and (w3932, x0_c, x2, x3_c, x4, x5, x6_c, x8_c, x11, x13, x14_c, x15_c, x16_c, x17, x18_c, x20, x21_c, x22_c, x24_c, x25_c, x26, x28_c, x29_c, x30_c, x34, x35_c, x36_c, x38, x41_c, x42_c, x43, x44_c, x47_c, x48_c, x50, x51, x52_c, x53_c, x54, x56, x57_c, x60, x61_c, x62_c, x63, x67, x68_c, x69_c, x70_c, x72_c, x73_c, x74_c, x76, x78, x79_c, x80, x84, x85, x86_c, x89_c, x91_c, x92, x93_c, x94, x95, x96_c, x98_c, x99_c);
and (w3933, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57_c, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3934, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3935, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79, x80);
and (w3936, x16_c, x26_c, x34_c, x45, x73_c, x75_c, x78_c, x79, x81, x83_c, x88, x91_c);
and (w3937, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x95_c, x97_c);
and (w3938, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3939, x0_c, x1, x2_c, x4, x5_c, x6_c, x8, x9_c, x10, x11, x12, x13, x16, x17, x18_c, x19, x21, x22_c, x23, x24_c, x25_c, x26, x30_c, x31, x32, x34_c, x35, x39, x42, x44, x46_c, x47_c, x48, x49_c, x51, x52_c, x53, x54, x56, x57_c, x58_c, x59_c, x61, x63, x64, x66, x67, x68, x72_c, x73, x74, x75, x77_c, x79, x80_c, x81, x82, x83, x84, x85_c, x86, x87_c, x88_c, x89_c, x90, x92, x94, x97, x98_c, x99_c);
and (w3940, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w3941, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x77_c, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3942, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3943, x0_c, x3_c, x4, x6_c, x10_c, x11, x13_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3944, x0_c, x1, x2, x3, x4, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3945, x14, x94);
and (w3946, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x85, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3947, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94, x95, x97_c);
and (w3948, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63, x75, x84_c, x85_c, x97_c);
and (w3949, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3950, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x40, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3951, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w3952, x4_c, x5, x6_c, x22, x31, x51_c, x59_c, x61, x64, x66, x70_c, x75_c, x79_c, x81_c, x82_c);
and (w3953, x12_c, x40, x42_c, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w3954, x4_c, x9_c, x11_c, x12, x25, x27, x50, x56, x58_c, x71, x81_c, x88_c, x93_c, x95_c);
and (w3955, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78, x84_c, x85_c, x97_c);
and (w3956, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3957, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x97, x98, x99_c);
and (w3958, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w3959, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89, x91_c, x92_c, x94, x95_c, x97_c);
and (w3960, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x38, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3961, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3962, x4_c, x5, x7_c, x12, x14, x15, x21_c, x23_c, x30_c, x31, x36_c, x37_c, x41_c, x45_c, x49, x51, x52, x54_c, x55, x61, x62_c, x66_c, x70, x75_c, x77_c, x90_c, x92, x96);
and (w3963, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3964, x4_c, x10, x15_c, x21, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w3965, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w3966, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x93_c, x95_c, x98, x99_c);
and (w3967, x11, x12_c, x15, x17_c, x23_c, x24, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3968, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33, x40, x82, x90_c, x96, x98, x99_c);
and (w3969, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x57, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w3970, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3971, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x88, x90_c, x91, x92, x95, x97_c);
and (w3972, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3973, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w3974, x0_c, x1_c, x2_c, x3_c, x4_c, x6, x7_c, x8_c, x9, x11, x12, x17, x19_c, x20_c, x21, x22, x24_c, x25_c, x27_c, x29_c, x30_c, x31_c, x32, x33, x37_c, x39, x42, x44, x45, x46_c, x49, x50, x51_c, x52_c, x53_c, x55, x57, x61_c, x63, x66, x67_c, x69_c, x70, x72, x73_c, x76, x77_c, x79, x80_c, x81, x83_c, x85_c, x87, x88_c, x90_c, x92, x96, x98_c);
and (w3975, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91, x92, x93_c, x94_c, x97_c);
and (w3976, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3977, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3978, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3979, x2_c, x11, x13_c, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3980, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x76_c, x85, x89, x93, x97_c, x98_c, x99_c);
and (w3981, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x49, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w3982, x2_c, x3, x5, x6, x7, x8, x9_c, x10_c, x12, x13, x14_c, x16_c, x21, x24_c, x27_c, x29_c, x30, x32, x34, x35, x38, x40, x42, x44_c, x45, x48, x49, x50_c, x51_c, x52, x53, x55, x56, x59, x61, x62, x63, x67_c, x68, x70, x74, x78, x83, x84_c, x86_c, x88_c, x89_c, x91, x96, x97, x98_c);
and (w3983, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x44_c, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w3984, x2_c, x4_c, x5, x6_c, x9, x10_c, x12_c, x16, x18, x19, x20_c, x21_c, x22, x24, x25_c, x26, x27_c, x28, x31, x32_c, x33, x34, x36, x37, x38_c, x39, x40_c, x41, x44, x45, x46_c, x47_c, x48, x49, x50, x51, x52, x53_c, x54, x56, x57_c, x58_c, x60, x61_c, x62, x64_c, x65_c, x66, x67_c, x70, x71, x72_c, x74, x76, x80, x81_c, x83, x85, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93, x98, x99);
and (w3985, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x97_c, x98, x99_c);
and (w3986, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w3987, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x85, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w3988, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22_c, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3989, x0, x3, x8, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w3990, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w3991, x1, x4, x5_c, x13_c, x15, x23, x24_c, x31, x33, x39_c, x43, x46, x49_c, x50_c, x54_c, x60_c, x67, x71_c, x74_c, x78_c, x83_c, x86_c, x87, x89_c, x93, x95_c);
and (w3992, x5_c, x9, x27, x51_c, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w3993, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3994, x2_c, x3, x4_c, x6_c, x7_c, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w3995, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x59_c, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w3996, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w3997, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w3998, x51_c, x58_c, x65);
and (w3999, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4000, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94, x95, x96, x97_c);
and (w4001, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62_c, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4002, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4003, x12_c, x32, x47_c, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4004, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x95_c, x96, x98, x99);
and (w4005, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x54, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4006, x0, x1, x3, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x13_c, x14, x15, x16_c, x17, x18_c, x20, x22_c, x23, x25_c, x29, x33_c, x35, x36_c, x38, x39_c, x41_c, x42, x43, x44, x45_c, x46, x47_c, x48_c, x54, x55, x58_c, x59, x60_c, x63, x68, x69_c, x70, x73_c, x74_c, x75_c, x76_c, x77, x79_c, x81, x82, x84_c, x92_c, x96_c, x98, x99_c);
and (w4007, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x57_c, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4008, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x22, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4009, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4010, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4011, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87_c, x89, x93, x97_c);
and (w4012, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x84_c, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4013, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4014, x5, x10, x16, x21_c, x32_c, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w4015, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x20, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4016, x0_c, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4017, x1_c, x6, x8, x10, x20, x24, x27_c, x28, x29, x34, x35, x40, x43_c, x44, x45_c, x46_c, x48_c, x49_c, x53, x59_c, x61, x63, x67_c, x69_c, x70, x71_c, x77, x79_c, x80, x91, x96_c);
and (w4018, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32_c, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4019, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x88, x90_c, x91, x92, x95, x97_c);
and (w4020, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4021, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4022, x13, x22, x36_c, x38, x42_c, x54_c, x60, x77, x84, x88_c, x89_c);
and (w4023, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x47_c, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4024, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4025, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43, x82, x90_c, x96, x98, x99_c);
and (w4026, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4027, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x58_c, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4028, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91_c, x93_c, x95_c, x96, x98, x99);
and (w4029, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4030, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4031, x11, x12_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4032, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x93_c, x96, x99_c);
and (w4033, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4034, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4035, x1, x4_c, x7, x8_c, x11_c, x14, x15_c, x17, x18_c, x21_c, x22, x24, x25_c, x28_c, x31, x32, x34, x35, x38_c, x39_c, x41_c, x42, x48_c, x49, x50, x52, x57, x61_c, x62_c, x63_c, x64_c, x66_c, x67_c, x68_c, x69_c, x71_c, x73_c, x76, x77, x78_c, x80_c, x81, x82_c, x83, x84_c, x87_c, x93_c, x94, x97_c, x99);
and (w4036, x7_c, x12_c, x17_c, x19, x36_c, x41, x59, x64, x84, x91, x98_c, x99_c);
and (w4037, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88, x93_c, x97_c);
and (w4038, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4039, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4040, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4041, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x65_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4042, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x88_c, x90, x93_c, x95_c, x96, x98, x99);
and (w4043, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4044, x12_c, x32, x89, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4045, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88, x89_c, x90, x91_c, x92_c, x93, x95_c, x96_c, x98, x99_c);
and (w4046, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x77_c, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4047, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x52, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w4048, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4049, x0_c, x1_c, x4, x6, x7, x8, x9_c, x10_c, x11_c, x15_c, x16, x18_c, x20, x21, x22_c, x23, x24, x25_c, x27, x28_c, x29, x30, x32, x34, x36_c, x37_c, x38_c, x39_c, x40_c, x41, x42, x43_c, x44, x46_c, x47, x48_c, x49, x50_c, x52_c, x54_c, x55_c, x56, x57, x59, x60, x62, x64, x65, x67, x68, x71_c, x72_c, x73, x74, x76, x77, x80, x81, x82, x83, x84, x87, x90_c, x91, x92, x93_c, x94, x95_c, x96, x97, x98, x99_c);
and (w4050, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4051, x4_c, x10, x15_c, x21, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4052, x2_c, x4, x5, x6_c, x11_c, x13, x16, x21, x23, x31, x32_c, x33_c, x34, x36, x38_c, x40, x43_c, x46_c, x47, x48_c, x50_c, x56_c, x61, x62_c, x65_c, x67, x68_c, x73_c, x74_c, x77_c, x78, x80_c, x82, x83, x85, x88_c, x89_c, x90_c, x92, x93, x95, x96_c, x97_c);
and (w4053, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4054, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4055, x0_c, x1_c, x2, x4, x5, x8, x9, x10_c, x11, x13, x14_c, x15_c, x17_c, x18, x20_c, x21, x22, x23_c, x26_c, x27, x28, x29_c, x30_c, x33, x35, x36, x37_c, x38, x39, x40_c, x41_c, x44, x45_c, x46, x49_c, x50_c, x52, x53_c, x54, x56_c, x57, x58, x60, x61_c, x62_c, x65_c, x66, x69, x72_c, x73, x74, x75_c, x79, x81_c, x85, x87, x88_c, x91_c, x93, x95_c, x96, x97_c, x98, x99_c);
and (w4056, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x69, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4057, x0, x1, x2, x3, x4, x5_c, x7_c, x8_c, x9_c, x10_c, x13, x14, x15_c, x16, x17, x18, x19_c, x23, x24, x25, x26_c, x27, x28, x29, x30, x31_c, x32_c, x33, x34_c, x36_c, x37, x39, x43_c, x44, x45_c, x46_c, x47, x48, x50_c, x51, x52, x53_c, x54_c, x55_c, x56_c, x58, x59_c, x62, x63_c, x64, x65, x67, x69_c, x70, x71_c, x73_c, x74, x75_c, x76, x79, x80_c, x81, x82, x84, x85, x86_c, x87_c, x92, x93, x94_c, x95, x97_c, x98, x99_c);
and (w4058, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4059, x1_c, x3_c, x7_c, x8, x9_c, x10_c, x11_c, x12, x16_c, x17, x18_c, x23_c, x25_c, x26_c, x27, x30_c, x31, x32_c, x33_c, x40, x42, x44_c, x45_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52, x55, x56_c, x57, x58_c, x61_c, x62_c, x65_c, x66_c, x69_c, x70, x72, x73_c, x75_c, x77, x79_c, x80_c, x81, x86, x88, x90, x91, x92_c, x96_c, x97_c, x99_c);
and (w4060, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60_c, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4061, x0_c, x5, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4062, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4063, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4064, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4065, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4066, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x92, x96_c, x98);
and (w4067, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4068, x2_c, x3, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4069, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x19, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4070, x0_c, x3_c, x6, x7, x10_c, x11_c, x12, x13, x15, x16_c, x18_c, x19_c, x23_c, x26, x34, x39, x40, x47_c, x49, x53, x54, x57_c, x61, x62_c, x63, x64_c, x66, x67, x69_c, x77, x78_c, x80_c, x81, x86, x87, x89_c, x90_c, x92, x94, x95, x98, x99);
and (w4071, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4072, x0, x2, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4073, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x23_c, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4074, x2_c, x11, x18_c, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4075, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x76, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4076, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w4077, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4078, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98_c);
and (w4079, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61, x83_c);
and (w4080, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4081, x12_c, x40, x82, x90_c, x92_c, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4082, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4083, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x63_c, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4084, x0, x1, x3, x4, x5_c, x6, x7_c, x8_c, x9_c, x10, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23, x24_c, x25, x26, x27_c, x28_c, x29_c, x30_c, x31_c, x32, x33, x34_c, x35, x36, x37_c, x38, x39_c, x40_c, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x50, x51_c, x52, x53, x54, x55_c, x56, x57_c, x58, x59, x60, x61, x62, x63, x64, x65_c, x66_c, x67, x68, x69, x70, x71, x72, x73, x74_c, x75, x76, x77_c, x78, x79, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92, x93, x94, x95, x96, x97_c, x98, x99_c);
and (w4085, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4086, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x79, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4087, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4088, x6, x17_c, x20, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w4089, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4090, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4091, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x90, x93, x94_c, x96, x97);
and (w4092, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78, x82, x83, x93_c, x97_c);
and (w4093, x36, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4094, x2_c, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4095, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4096, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93_c, x95, x96, x97, x99_c);
and (w4097, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x59, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4098, x2, x9_c, x14, x21, x29_c, x36_c, x50, x70_c, x93, x96_c);
and (w4099, x0_c, x1, x2_c, x3_c, x4_c, x5_c, x6, x7_c, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16, x17_c, x18, x19_c, x20, x21, x22_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x35, x36_c, x37, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46_c, x47, x48, x49_c, x50_c, x51, x52_c, x53, x54_c, x55, x56_c, x57, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65_c, x66_c, x67, x68, x69_c, x70_c, x71_c, x72, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80, x81_c, x82, x83_c, x84_c, x85, x86_c, x87_c, x88, x89, x91, x92_c, x93_c, x94_c, x95_c, x96_c, x98_c, x99_c);
and (w4100, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24_c, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4101, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4102, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4103, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4104, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x79_c, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4105, x6, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4106, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75, x83_c);
and (w4107, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70_c, x83_c);
and (w4108, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25_c, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4109, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31_c, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4110, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69, x72_c, x81, x84, x85, x95, x99);
and (w4111, x0, x4_c, x10, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4112, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x90_c, x91_c, x93_c, x95_c, x96, x98, x99);
and (w4113, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4114, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75_c, x81, x84, x85, x95, x99);
and (w4115, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x75, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4116, x12_c, x20, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4117, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4118, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4119, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x38, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4120, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85, x90_c, x93_c, x97_c);
and (w4121, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4122, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4123, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92, x93_c, x95_c, x96_c, x97_c);
and (w4124, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x61_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4125, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x65_c, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4126, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x87, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4127, x0, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4128, x24_c, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4129, x5_c, x9, x25, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4130, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4131, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x42, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4132, x0, x1, x2_c, x3, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w4133, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4134, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4135, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4136, x12_c, x19, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4137, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x36, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4138, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x47, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4139, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x23, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4140, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78_c, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4141, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x51_c, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4142, x0, x1, x3_c, x4, x7, x8_c, x9_c, x10_c, x11, x12_c, x14_c, x15_c, x16_c, x17_c, x18, x19, x21, x22_c, x25_c, x27_c, x29, x30_c, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x45_c, x46_c, x47_c, x48, x49, x50, x52, x53_c, x55, x56_c, x57, x58_c, x59, x60_c, x61, x62, x64, x65, x66, x67, x68_c, x70_c, x72, x73_c, x74_c, x75, x76_c, x77, x78_c, x79, x80_c, x81_c, x82_c, x83, x84_c, x85, x86_c, x87, x89, x90, x91, x93, x95_c, x96_c, x97_c, x98, x99);
and (w4143, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45_c, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w4144, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4145, x1, x2_c, x6, x7_c, x9, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4146, x0_c, x1_c, x2_c, x3_c, x4_c, x6, x7_c, x8_c, x9, x10, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21_c, x22, x23, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45_c, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x55_c, x56, x57_c, x58, x59, x60_c, x61, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75_c, x76, x77, x78, x79, x80_c, x81_c, x82, x83_c, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95_c, x96, x97_c, x98_c, x99_c);
and (w4147, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69, x71_c);
and (w4148, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4149, x12_c, x14, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4150, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4151, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x71, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4152, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x84, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4153, x0_c, x5_c, x9, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4154, x8, x21, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4155, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4156, x11_c, x15_c, x16, x18, x21, x28_c, x35, x71_c);
and (w4157, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42, x82, x90_c, x96, x98, x99_c);
and (w4158, x2_c, x11, x25, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4159, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x50_c, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4160, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4161, x0_c, x6, x10, x17_c, x29_c, x52, x58_c, x74_c, x89, x92_c, x96, x97);
and (w4162, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4163, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x41, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4164, x28_c, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4165, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29, x83_c);
and (w4166, x3, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w4167, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4168, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x93, x97_c);
and (w4169, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x91_c, x95_c, x96, x98, x99);
and (w4170, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x65_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4171, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4172, x12_c, x40, x58_c, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4173, x5_c, x9, x27, x44_c, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4174, x1, x2, x3, x7, x8_c, x9_c, x10_c, x11, x13, x15, x16, x18_c, x21, x22_c, x23, x26_c, x27_c, x29_c, x31, x32_c, x34, x37, x38, x39_c, x40, x41_c, x42_c, x43, x45, x49_c, x50_c, x51, x53, x56, x57, x58_c, x61_c, x62_c, x63, x64_c, x68_c, x69, x70, x72, x75_c, x76, x77, x79, x81_c, x84, x87, x92_c, x95, x97, x98_c);
and (w4175, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96_c);
and (w4176, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x63, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4177, x4_c, x5_c, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w4178, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4179, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83_c, x90_c, x93_c, x97_c);
and (w4180, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4181, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4182, x2, x3_c, x4_c, x15, x24, x34, x36_c, x39_c, x41_c, x42_c, x47, x52, x54, x56_c, x57, x68, x69_c, x70, x81, x82, x86_c, x92, x97_c, x99);
and (w4183, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4184, x12_c, x17, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4185, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4186, x11, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4187, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4188, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4189, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x64, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4190, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4191, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4192, x6, x13, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4193, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x31, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4194, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89_c, x93_c, x97_c);
and (w4195, x1_c, x3_c, x4, x10_c, x12_c, x13_c, x15_c, x36, x38_c, x39, x42_c, x43_c, x48, x52_c, x57, x58_c, x59, x60_c, x63, x65_c, x68_c, x76, x82, x86_c, x99_c);
and (w4196, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x96_c, x98, x99);
and (w4197, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49_c, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4198, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x96, x97_c, x98_c, x99_c);
and (w4199, x0_c, x2_c, x3, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4200, x11_c, x15_c, x16_c, x23_c, x71_c);
and (w4201, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42, x83_c);
and (w4202, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x80_c, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4203, x40, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4204, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x84_c, x85_c, x96_c, x98, x99_c);
and (w4205, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37_c, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4206, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4207, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4208, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4209, x0_c, x5, x12, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4210, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4211, x0, x4_c, x12_c, x22_c, x27_c, x30, x32_c, x39, x43_c, x48, x54, x69_c, x78_c, x92, x96);
and (w4212, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x83, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4213, x12_c, x32, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4214, x0, x3, x10, x13, x14, x15, x16_c, x22, x35, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4215, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x87_c, x89, x90_c, x91, x93, x94_c, x95_c, x96, x97);
and (w4216, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x35, x36, x37, x38_c, x39_c, x40_c, x41_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4217, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x40, x82, x90_c, x96, x98, x99_c);
and (w4218, x13_c, x15, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w4219, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57, x73_c, x76, x85, x89, x93, x97_c);
and (w4220, x0, x2, x4, x5_c, x6, x8, x9_c, x12, x13, x15_c, x16, x17_c, x18_c, x19, x22_c, x23_c, x25_c, x27_c, x28, x29_c, x30_c, x31_c, x33_c, x35_c, x36, x38, x40, x41, x42_c, x43_c, x45_c, x46, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x56_c, x58, x61_c, x62, x63, x65, x68, x69_c, x70, x71_c, x73, x75, x76_c, x78_c, x79_c, x80, x82_c, x83_c, x86_c, x90, x91, x92_c, x93, x94_c, x96, x97);
and (w4221, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4222, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x81, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4223, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4224, x2, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4225, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4226, x0, x1, x2, x3_c, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4227, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4228, x2, x3, x4, x6_c, x7_c, x8, x9, x10, x12_c, x16, x17_c, x18_c, x20_c, x21, x22_c, x24_c, x25, x27_c, x28_c, x29_c, x30_c, x32, x34_c, x35_c, x36, x38_c, x40_c, x41, x44_c, x45, x46, x47_c, x50, x51_c, x52_c, x55_c, x56_c, x57, x58, x60, x61_c, x65_c, x66, x67_c, x68_c, x69_c, x70_c, x72, x75, x76, x77_c, x78_c, x79, x80, x81, x82_c, x85_c, x86_c, x87, x88_c, x89, x91, x92_c, x94_c, x95_c, x96, x97_c, x98_c);
and (w4229, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4230, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4231, x0, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x8, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18, x19, x20, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34_c, x35, x36, x37_c, x38_c, x39, x40_c, x41, x42_c, x43, x44, x45, x46_c, x47_c, x48, x49, x50, x51_c, x52_c, x53_c, x54, x55_c, x56_c, x57, x58_c, x59, x60, x61_c, x62_c, x63, x64, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81, x82, x83, x84_c, x85_c, x86_c, x87, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w4232, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87_c, x97_c);
and (w4233, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4234, x0_c, x1, x2, x4, x14, x16, x17_c, x20_c, x22_c, x23_c, x25, x31_c, x33_c, x38_c, x44, x45_c, x47, x53, x54_c, x55, x56_c, x57_c, x61_c, x63_c, x70_c, x74, x78_c, x83_c, x84, x85_c, x86, x90_c, x92_c, x94_c, x95, x96, x97, x99);
and (w4235, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4236, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x70, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4237, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4238, x1_c, x2_c, x4_c, x5, x7_c, x8_c, x9_c, x10_c, x14, x15_c, x16, x17_c, x18_c, x20_c, x23, x25, x26_c, x28_c, x30, x31_c, x32, x37, x38, x44, x45_c, x47, x48, x52_c, x53, x54, x55, x57, x58, x59, x65, x66_c, x67_c, x68_c, x69_c, x71_c, x72, x73, x77, x79, x80, x81_c, x84, x85_c, x86, x87_c, x88, x90_c, x91_c, x92_c, x93, x96, x98, x99_c);
and (w4239, x0_c, x5_c, x6, x12_c, x16, x17_c, x18_c, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4240, x0_c, x1, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4241, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4242, x7, x16_c, x21, x24, x26, x37_c, x40, x41_c, x44, x48_c, x53, x64_c, x74, x76_c, x78_c, x80, x82_c, x86_c, x90_c, x91, x94_c, x95);
and (w4243, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x74_c, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4244, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4245, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4246, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4247, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4248, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4249, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x67_c, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w4250, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52_c, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4251, x0, x2, x5_c, x6, x7_c, x8, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4252, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15, x16, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4253, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x91_c, x93, x95_c, x96_c, x98_c);
and (w4254, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4255, x5, x10, x16_c, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w4256, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4257, x2, x5, x6_c, x8_c, x9_c, x13_c, x14_c, x15_c, x16, x17, x18_c, x22, x23_c, x24_c, x28_c, x29, x30_c, x31_c, x34, x35, x36_c, x37, x38_c, x39, x40_c, x41_c, x42, x44_c, x45_c, x46_c, x47_c, x49, x51_c, x54, x55_c, x56_c, x57, x58, x59_c, x60_c, x62_c, x64, x65_c, x66_c, x69, x72_c, x74, x75_c, x79, x80_c, x82, x83, x85, x87, x88, x89, x90_c, x92, x93_c, x95, x97_c, x98, x99);
and (w4258, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x66_c, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4259, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x98, x99);
and (w4260, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4261, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4262, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70_c, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4263, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4264, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4265, x1, x6, x7_c, x12_c, x13, x22_c, x23_c, x25_c, x27, x28_c, x31, x32_c, x33_c, x37_c, x39_c, x40_c, x43, x44, x49, x55_c, x58_c, x61, x63_c, x64_c, x67_c, x68, x70, x75, x78_c, x88, x89_c, x90, x91_c, x94, x98);
and (w4266, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x83_c, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4267, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4268, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4269, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4270, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x10, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4271, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4272, x0, x1_c, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4273, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4274, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x33_c, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4275, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x61_c, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4276, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4277, x1, x2_c, x6, x7_c, x8, x10, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4278, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4279, x4_c, x10, x15_c, x20_c, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w4280, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x49, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4281, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4282, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x19, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w4283, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4284, x12_c, x32, x50_c, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4285, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4286, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x91_c, x92, x95, x97_c);
and (w4287, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x47_c, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4288, x0_c, x1, x2, x3_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4289, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25, x83_c);
and (w4290, x4_c, x10, x15_c, x22_c, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w4291, x1_c, x2, x3, x4, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4292, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4293, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4294, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4295, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x60_c, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4296, x1, x3_c, x4_c, x5_c, x6_c, x7, x9, x10_c, x11, x12_c, x13, x15, x17_c, x18_c, x19, x21, x23_c, x24_c, x25_c, x26, x27, x28, x29, x33_c, x34, x35, x36_c, x37_c, x39, x41_c, x42, x43, x44_c, x45, x49, x51, x52_c, x53, x54_c, x55, x57_c, x59_c, x60, x61_c, x63_c, x64_c, x65, x67_c, x69, x70_c, x71, x73, x75_c, x77, x78, x79_c, x80_c, x81, x82_c, x83, x87, x88_c, x89_c, x91_c, x92_c, x93, x94, x95, x96_c, x98, x99);
and (w4297, x8, x21_c, x25_c, x27_c, x30_c, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4298, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4299, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81, x85, x89, x93, x97_c);
and (w4300, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4301, x0_c, x1_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4302, x0_c, x1, x2_c, x3, x4_c, x6, x7, x8_c, x12_c, x13, x14_c, x15, x16, x17, x20, x21_c, x23_c, x24, x25, x26, x27_c, x28_c, x30_c, x31_c, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x40, x42, x43_c, x44, x45_c, x46_c, x49_c, x50_c, x51_c, x52, x53, x54, x55_c, x57, x58_c, x63, x64, x65_c, x66_c, x67, x69, x71, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79_c, x84_c, x88_c, x90, x91, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4303, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33, x83_c);
and (w4304, x4_c, x10, x15_c, x16, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w4305, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4306, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x32, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4307, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4308, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4309, x0_c, x3_c, x4_c, x6, x7, x10_c, x11, x13_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4310, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x27, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4311, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4312, x2_c, x4, x5, x7_c, x9_c, x13_c, x14_c, x18_c, x19, x20_c, x22_c, x24_c, x28_c, x30, x32, x35_c, x36_c, x37_c, x38, x40, x44, x47_c, x48, x50, x52_c, x59, x61_c, x63_c, x65, x71_c, x72, x73, x76_c, x77, x79_c, x80, x81, x83, x84, x87_c, x89_c, x93, x94_c, x97, x98);
and (w4313, x2, x6, x7, x12_c, x14_c, x29_c, x31, x32, x33_c, x34_c, x35, x36, x37_c, x40, x41_c, x43, x44, x45, x46_c, x47, x53_c, x55, x56_c, x65, x74, x75, x76_c, x78, x81_c, x82, x83_c, x86, x87, x88_c, x90, x91, x92_c, x95_c, x97);
and (w4314, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4315, x0_c, x4_c, x5_c, x6, x12_c, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4316, x0, x1_c, x2, x4_c, x5_c, x6, x7, x8, x9, x11, x12, x13_c, x14, x16, x17, x18, x19_c, x21, x22_c, x23_c, x24_c, x25, x26, x27_c, x28_c, x29, x30_c, x31_c, x32, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40, x41_c, x43, x44, x45, x47_c, x48_c, x49, x50_c, x51_c, x52, x54, x56, x57, x58_c, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66, x67, x68, x69, x70, x73_c, x74, x75, x76_c, x77_c, x78, x79_c, x80, x81_c, x82, x84_c, x85, x86_c, x87, x88_c, x90, x91, x92_c, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w4317, x0, x1_c, x4_c, x7, x17_c, x18_c, x52_c, x66_c, x67_c, x70_c, x74_c, x99_c);
and (w4318, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4319, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4320, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x76, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4321, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87_c, x90_c, x91, x92, x95, x97_c);
and (w4322, x6, x13, x18, x20, x22_c, x31, x34_c, x38, x44_c, x46_c, x47_c, x54, x58, x61, x64, x68_c, x71_c, x74_c, x75_c, x76_c, x79, x80, x81, x99);
and (w4323, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4324, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x99);
and (w4325, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4326, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x40_c, x82, x90_c, x96, x98, x99_c);
and (w4327, x0, x1, x2, x5, x6_c, x7_c, x9_c, x11, x13_c, x14_c, x17, x18_c, x19_c, x20, x21, x22, x27_c, x29_c, x32, x33, x36, x38, x40, x41, x42_c, x43_c, x45_c, x46, x49_c, x50_c, x51_c, x52_c, x55_c, x57, x58_c, x60_c, x61_c, x63_c, x64, x65_c, x67, x69_c, x72_c, x74, x75_c, x77, x78, x79_c, x80, x81, x82, x83_c, x86_c, x90, x91_c, x92, x94_c, x96_c, x97, x99_c);
and (w4328, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4329, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w4330, x8, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4331, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x91_c, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4332, x12_c, x40, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4333, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4334, x0_c, x5, x23_c, x30, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4335, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x65, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4336, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80_c, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w4337, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4338, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48_c, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w4339, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x82_c, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4340, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4341, x3, x13, x24, x27_c, x29, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4342, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18_c, x40, x82, x90_c, x96, x98, x99_c);
and (w4343, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4344, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x73_c, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4345, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4346, x0, x2_c, x3, x5_c, x6, x9, x14_c, x15, x16, x18_c, x19, x20_c, x24, x26, x27, x28_c, x31, x39, x43, x47, x48, x50, x51, x65, x68_c, x69_c, x71_c, x72_c, x73, x74_c, x79, x80_c, x81, x86_c, x87, x96, x97, x99);
and (w4347, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48_c, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w4348, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30_c, x40, x82, x90_c, x96, x98, x99_c);
and (w4349, x3_c, x5, x6, x7_c, x10, x11, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4350, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4351, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x74, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4352, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4353, x5, x10, x16, x21_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4354, x3_c, x4, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4355, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4356, x0_c, x2_c, x6_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w4357, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4358, x8, x17, x18_c, x27_c, x34, x39_c, x55, x56_c, x61_c, x62_c, x70_c, x88_c);
and (w4359, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75_c, x82, x90_c, x96, x98, x99_c);
and (w4360, x0, x1, x2, x3, x4, x5_c, x6_c, x7, x8_c, x9, x10_c, x11, x12, x13_c, x14_c, x15_c, x17_c, x24, x25, x26_c, x29_c, x30_c, x31, x32_c, x33, x34_c, x35, x36, x37, x38_c, x41, x42_c, x43, x44_c, x46_c, x47_c, x48_c, x49_c, x50_c, x53, x54_c, x55, x57_c, x58, x59_c, x61, x62, x63_c, x64_c, x65_c, x68, x71_c, x72_c, x74_c, x75, x76, x79_c, x80, x81, x82_c, x84, x90, x94_c, x98);
and (w4361, x0, x3, x4, x8_c, x11_c, x12, x13_c, x14, x17_c, x18_c, x19, x22_c, x23_c, x26_c, x27, x28, x29_c, x30, x31, x33, x34_c, x36_c, x37, x38, x40, x43_c, x45_c, x47_c, x48_c, x49, x50_c, x51_c, x52, x53_c, x57, x58_c, x60, x64, x68, x71_c, x74_c, x75, x78_c, x79_c, x80, x83_c, x84, x86_c, x89_c, x92, x93_c, x94_c, x95_c);
and (w4362, x3_c, x9, x10_c, x13, x16, x17, x19, x20, x21, x25_c, x28, x30, x34_c, x35, x39, x41_c, x44_c, x46_c, x48, x50, x54, x55, x60_c, x61_c, x62_c, x63, x65, x67_c, x68_c, x70, x71_c, x73, x75, x78, x79_c, x81_c, x82, x83_c, x87_c, x89_c, x93_c, x97_c);
and (w4363, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4364, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x22_c, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4365, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4366, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4367, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4368, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4369, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4370, x8, x21_c, x25_c, x27_c, x34, x39_c, x42_c, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4371, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x66_c, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4372, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4373, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4374, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4375, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x15, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4376, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x51, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4377, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x80, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w4378, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4379, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x40, x82, x90_c, x96, x98, x99_c);
and (w4380, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4381, x0_c, x1, x2, x3_c, x4_c, x5_c, x6, x7, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15, x16_c, x17, x18, x19_c, x20, x21_c, x22_c, x23, x24, x25, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x42_c, x43, x45_c, x46_c, x47, x48_c, x50_c, x51, x52_c, x53_c, x54, x55, x56_c, x57_c, x58_c, x59_c, x60, x61, x62_c, x63_c, x64, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x72, x73, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81_c, x82, x83, x84, x85, x86, x87_c, x88, x90_c, x91, x92_c, x93_c, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w4382, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x95_c, x96_c, x98, x99);
and (w4383, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x34_c, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w4384, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x93, x95_c, x96, x98, x99);
and (w4385, x1_c, x4, x13, x17, x20, x29_c, x32, x37, x60, x65, x67_c, x69_c, x75, x76_c, x84_c, x91_c, x94);
and (w4386, x12_c, x18_c, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4387, x0, x1, x2_c, x3, x4_c, x5, x6, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15, x16, x17, x18, x19, x20, x21, x22_c, x23_c, x24, x25, x26_c, x27_c, x28, x29_c, x30_c, x31_c, x32, x33, x34, x35_c, x36, x37_c, x38_c, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x51, x52_c, x53, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61, x62_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69, x70, x71_c, x72, x73_c, x74_c, x75, x76, x77_c, x78, x79_c, x80, x81_c, x82, x83_c, x85, x86_c, x87_c, x88_c, x89, x90, x91, x92_c, x93_c, x94_c, x95_c, x96, x97, x98_c, x99_c);
and (w4388, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4389, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4390, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x76_c, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4391, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4392, x49, x80, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4393, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x88_c, x89, x91, x93_c, x94_c, x96, x97, x98, x99);
and (w4394, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x59_c, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4395, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x48, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4396, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4397, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4398, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x90_c, x93_c, x95_c, x96, x97_c, x98, x99);
and (w4399, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4400, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x88_c, x89, x91, x92, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4401, x0, x2_c, x3_c, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4402, x2, x3_c, x4_c, x5_c, x7_c, x8_c, x9, x10, x11, x12, x13_c, x14, x15_c, x16, x17_c, x18, x19_c, x20_c, x24_c, x25, x26_c, x27_c, x28_c, x29, x30, x31, x33_c, x34_c, x35, x36_c, x37_c, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45, x46, x47, x49, x50_c, x52, x54_c, x55_c, x56, x57_c, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x78_c, x79, x80_c, x82, x85_c, x86, x87, x88_c, x89_c, x90_c, x93_c, x94_c, x95, x96, x97, x98_c, x99_c);
and (w4403, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4404, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4405, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4406, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86, x93_c, x97_c);
and (w4407, x0, x1, x2_c, x4_c, x5, x6, x7_c, x9_c, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x18, x19, x20, x22_c, x23, x25, x27, x28, x29_c, x30_c, x31, x32, x33_c, x34_c, x35_c, x37, x39, x40, x41_c, x42_c, x43, x44_c, x45_c, x46, x47_c, x48_c, x50, x51_c, x52, x53, x54, x55_c, x56, x57_c, x58_c, x59, x60, x61_c, x62_c, x64, x65_c, x66_c, x70, x71_c, x73, x75_c, x77_c, x78_c, x79, x81, x82_c, x83_c, x89, x90_c, x91_c, x93, x95, x96_c, x97, x99);
and (w4408, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4409, x12_c, x40, x82, x90_c, x94, x95, x96_c, x98, x99_c);
and (w4410, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4411, x0_c, x1, x2_c, x3_c, x4, x5_c, x6, x7_c, x9_c, x10, x11, x12_c, x13_c, x14, x15_c, x16_c, x17, x18_c, x19_c, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x29, x30, x31, x32, x33, x34_c, x35_c, x36_c, x37, x38_c, x39_c, x40, x41, x42_c, x43, x44, x46_c, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54_c, x55, x57_c, x58_c, x59_c, x60, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x69_c, x70, x71, x72, x73_c, x74, x75_c, x76, x77, x78, x79, x80, x81_c, x82, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91_c, x92_c, x93, x94_c, x95_c, x97, x99_c);
and (w4412, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x52, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4413, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4414, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x16_c, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4415, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x95, x96_c, x97_c, x98, x99_c);
and (w4416, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x53, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4417, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w4418, x0, x2, x3, x6_c, x10_c, x11, x13_c, x19_c, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4419, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4420, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69_c, x73_c, x76, x85, x89, x93, x97_c);
and (w4421, x7_c, x12_c, x13, x25, x27, x31_c, x48_c, x49_c, x58, x59, x61_c, x62, x72_c, x73_c, x84_c, x87, x89_c, x90_c, x91_c);
and (w4422, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x50_c, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4423, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x73_c, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4424, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4425, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4426, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4427, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x89_c, x91_c, x92, x93, x94, x95, x96_c, x97_c);
and (w4428, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x20, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4429, x0, x3, x10, x13, x14, x15, x16_c, x22, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4430, x4_c, x5_c, x6_c, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4431, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x82_c, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4432, x0, x1_c, x2_c, x5_c, x6_c, x8, x16, x18, x24, x26_c, x28_c, x32, x35_c, x36, x38, x44, x45_c, x49_c, x50_c, x51, x56_c, x59_c, x62_c, x64_c, x65_c, x72, x73_c, x77, x80_c, x81_c, x82, x85_c, x87, x91_c, x92, x95_c, x96_c);
and (w4433, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91, x92, x93_c, x94, x96, x98_c, x99_c);
and (w4434, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79, x82, x83, x93_c, x97_c);
and (w4435, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x50_c, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w4436, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x66, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4437, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x93_c, x95_c, x96_c, x97, x98, x99_c);
and (w4438, x0_c, x2, x3_c, x4, x6_c, x7, x9, x10, x14_c, x15, x17, x18, x29_c, x31_c, x32, x33_c, x34, x35, x40_c, x43_c, x44, x46_c, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x56_c, x57, x58, x59_c, x60, x61_c, x62_c, x63, x64, x65_c, x66_c, x67, x68, x69_c, x70, x71_c, x72, x74, x76, x77_c, x78_c, x80, x81_c, x82, x83, x84_c, x85_c, x86, x87, x88, x89, x90_c, x92, x94, x95_c, x96_c, x99);
and (w4439, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4440, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x41_c, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4441, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4442, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w4443, x9_c, x14_c, x17, x24_c, x26_c, x56, x61, x73, x79);
and (w4444, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4445, x1_c, x2, x4, x5_c, x6_c, x8, x11, x12_c, x15, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4446, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4447, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4448, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w4449, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4450, x2_c, x3_c, x4_c, x6, x7, x8, x10_c, x12, x13, x16, x17_c, x18, x20_c, x21_c, x25_c, x26, x28_c, x36_c, x38_c, x39, x40, x41_c, x42_c, x43, x45, x46, x47_c, x61_c, x66, x70_c, x74_c, x76, x80, x81_c, x82_c, x83_c, x84_c, x87, x88_c, x90, x94_c, x97_c, x98);
and (w4451, x0, x1_c, x2, x3, x4_c, x6_c, x7, x8, x10, x11, x12, x13, x14, x15, x16_c, x17, x19_c, x20, x21_c, x22, x23_c, x24, x25, x27, x28_c, x29, x30_c, x31_c, x32, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40, x41_c, x42, x43_c, x44, x46_c, x47, x48_c, x49_c, x50, x51, x52_c, x53, x54_c, x55_c, x57, x58_c, x59, x60, x61_c, x62, x63, x64_c, x65, x66, x67_c, x68, x69, x70, x71, x72, x73, x74_c, x76_c, x77, x78_c, x79_c, x80, x81, x82_c, x83, x84, x85_c, x87_c, x88, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x98, x99_c);
and (w4452, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89, x90_c, x94_c, x95, x96_c, x97);
and (w4453, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4454, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4455, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87_c, x89, x93, x97_c);
and (w4456, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4457, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4458, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x89, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4459, x21_c, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4460, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4461, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34_c, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4462, x30_c, x64);
and (w4463, x0, x1, x3, x4_c, x5_c, x6, x8_c, x10_c, x12_c, x13, x15, x16, x20_c, x21, x23, x27_c, x28_c, x29_c, x30_c, x32_c, x33_c, x34_c, x36_c, x37_c, x44_c, x45, x47_c, x48_c, x49_c, x52, x53, x55_c, x56_c, x57, x58, x59, x61, x63_c, x65, x68, x69, x70, x71_c, x72, x73, x76, x79_c, x80, x81_c, x82, x84, x87_c, x89, x93_c, x96, x97_c, x98);
and (w4464, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x17, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4465, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4466, x40, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4467, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4468, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44_c, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4469, x5, x10, x16, x21_c, x30, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4470, x2_c, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4471, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x31_c, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4472, x12_c, x40, x52, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4473, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x77, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4474, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42_c, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4475, x0_c, x1_c, x2_c, x3_c, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12_c, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28_c, x29, x30_c, x31, x32, x33, x35_c, x36, x37_c, x38, x39, x41, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x52_c, x54, x55, x56, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x66, x67, x68, x69_c, x70_c, x71, x72, x74_c, x75, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87, x88_c, x89, x90, x91_c, x92, x93, x94, x97_c, x98_c, x99);
and (w4476, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x51, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4477, x7, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4478, x38, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4479, x12_c, x15, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4480, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4481, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4482, x0_c, x2_c, x4_c, x7_c, x9_c, x11_c, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4483, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4484, x69_c, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4485, x43, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4486, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w4487, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70, x75, x84_c, x85_c, x97_c);
and (w4488, x0, x2_c, x3, x4_c, x5_c, x6_c, x7, x10_c, x11, x12, x13, x14, x17, x18_c, x20_c, x21_c, x22_c, x24, x25_c, x26_c, x27, x28_c, x31_c, x32, x34, x35, x38, x39, x41, x44_c, x45_c, x46, x47, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58, x59, x60_c, x61, x62, x63, x64_c, x65_c, x66_c, x67, x68_c, x69, x71_c, x73, x75, x77, x78, x79_c, x80, x81, x83_c, x84_c, x85_c, x86_c, x88, x90_c, x91_c, x92_c, x93_c, x95, x98_c);
and (w4489, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x78_c, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4490, x2_c, x11, x29_c, x99_c);
and (w4491, x15, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4492, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x69_c, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4493, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4494, x0_c, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w4495, x13_c, x49, x64, x71, x72_c, x79_c, x81_c, x87, x90, x93_c, x97_c);
and (w4496, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x36_c, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4497, x5_c, x9, x27, x48_c, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4498, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x97_c, x98, x99_c);
and (w4499, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x89, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4500, x0, x3, x7, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4501, x0, x3, x5_c, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4502, x0_c, x3_c, x4_c, x6, x7_c, x10_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4503, x0_c, x4_c, x7_c, x9, x14_c, x20, x22_c, x23, x24_c, x27, x30_c, x31, x36_c, x39, x40, x43, x45, x46, x47_c, x51_c, x52_c, x53_c, x57, x58, x66_c, x69_c, x70, x71, x72_c, x73_c, x78, x83, x84_c, x86, x88, x90, x93, x94, x96_c, x97, x98);
and (w4504, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75_c, x76, x85, x89, x93, x97_c);
and (w4505, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45_c, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4506, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4507, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x41_c, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4508, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x22, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4509, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4510, x0_c, x5, x23_c, x30_c, x31, x32, x34_c, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4511, x0, x1_c, x2_c, x3_c, x4, x7_c, x10, x11_c, x12, x13, x14_c, x15, x16_c, x18_c, x20_c, x21_c, x22_c, x23, x24, x25_c, x26_c, x27, x28_c, x29, x30, x31_c, x32, x33, x34, x35, x36, x37_c, x38_c, x39_c, x40, x41, x42_c, x43_c, x45, x46, x47, x48, x49_c, x50, x51_c, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60, x61_c, x62, x63, x65, x66_c, x67_c, x68_c, x69, x71, x72_c, x73, x75, x76, x77, x78, x79, x80, x81_c, x82_c, x83, x84_c, x85_c, x86, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94, x95, x96_c, x97_c, x98, x99);
and (w4512, x0, x1, x2_c, x3_c, x4_c, x5, x6_c, x8_c, x10_c, x11, x12, x13, x14, x15_c, x16, x18_c, x19_c, x20, x21_c, x22_c, x26_c, x27_c, x28_c, x29_c, x31, x32, x33, x34_c, x36, x37_c, x38_c, x39_c, x40, x41, x42, x43, x44, x46_c, x47, x49, x50_c, x52_c, x53, x54, x55_c, x56_c, x57_c, x58, x59_c, x61_c, x62_c, x63, x64_c, x66_c, x67_c, x68_c, x73, x75_c, x76, x77_c, x78_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x86_c, x87_c, x88_c, x89, x90, x91_c, x92, x96_c, x97, x98_c);
and (w4513, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x17, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4514, x0_c, x2_c, x3_c, x4_c, x5_c, x6, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4515, x8, x21_c, x25_c, x27_c, x33_c, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4516, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w4517, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93_c);
and (w4518, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c, x99);
and (w4519, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4520, x12_c, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4521, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4522, x12_c, x32, x91, x92_c, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4523, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92, x93_c, x95_c);
and (w4524, x14, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4525, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4526, x6, x7_c, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4527, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x62, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4528, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4529, x0, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4530, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4531, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x20, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4532, x0, x1_c, x2_c, x3, x4_c, x6_c, x7_c, x8, x10, x11_c, x12_c, x13, x14, x15, x16, x17_c, x20_c, x22, x23_c, x25_c, x26_c, x27, x28, x29, x30_c, x31_c, x33_c, x34, x36, x37_c, x39_c, x40_c, x42_c, x43, x46, x47_c, x48_c, x49, x50, x51_c, x52_c, x53, x54, x55_c, x56, x57_c, x58_c, x59, x61_c, x62, x63_c, x64, x65_c, x68_c, x69_c, x71_c, x72_c, x73, x74_c, x75_c, x77, x78_c, x79_c, x82_c, x83_c, x84_c, x85, x87, x88_c, x89, x91_c, x92_c, x93, x94, x95, x96_c, x97_c, x98, x99_c);
and (w4533, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x66_c, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4534, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4535, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x90, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4536, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w4537, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x79_c, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4538, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x71, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4539, x5_c, x9, x23, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4540, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x90_c, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4541, x1_c, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4542, x2_c, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4543, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4544, x1_c, x2, x4, x5_c, x6, x11, x12_c, x15, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4545, x2_c, x11, x29_c, x48_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4546, x2_c, x3_c, x5, x7, x8_c, x9, x10_c, x11_c, x12_c, x13, x14_c, x16_c, x21_c, x23, x24_c, x25, x26_c, x28_c, x29, x30, x31_c, x32, x33, x34, x35_c, x37_c, x38, x39_c, x40_c, x41, x42, x43, x44_c, x45, x46_c, x47_c, x48_c, x51_c, x53_c, x54, x56, x57_c, x58_c, x59, x60, x61, x62_c, x63_c, x66_c, x68_c, x69, x70, x71_c, x72_c, x73, x74, x75, x76, x77_c, x79_c, x80, x81, x83_c, x84, x86_c, x87_c, x89, x90_c, x91, x92_c, x93_c, x95, x97, x98_c, x99_c);
and (w4547, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4548, x0_c, x1, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4549, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x82, x90_c, x96, x98, x99_c);
and (w4550, x9, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4551, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x58, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4552, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x81, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4553, x12_c, x32_c, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4554, x12_c, x32, x87, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4555, x0, x1, x2_c, x3, x4, x5, x6_c, x7, x9, x10_c, x11_c, x12_c, x13_c, x14, x15, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23, x24, x25, x26_c, x27, x28_c, x29_c, x30, x31, x32, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40, x41, x42_c, x43_c, x44, x45, x46, x47_c, x48, x49, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67, x68, x69_c, x70_c, x71, x72, x73, x74, x75, x76_c, x77, x79_c, x80_c, x81_c, x83_c, x84_c, x85, x87, x88, x89_c, x90_c, x91_c, x92_c, x93, x94, x95_c, x96_c, x97, x98_c, x99);
and (w4556, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4557, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4558, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x73, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4559, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4560, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4561, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4562, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4563, x3, x13, x23, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4564, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x50_c, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4565, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x60_c, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4566, x12_c, x22_c, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4567, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4568, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
assign w4569 = x2_c;
and (w4570, x0_c, x2_c, x4_c, x7, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4571, x0, x1, x2_c, x3_c, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w4572, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x40, x82, x90_c, x96, x98, x99_c);
and (w4573, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4574, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85, x93_c, x97_c);
and (w4575, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4576, x0_c, x1_c, x2_c, x3_c, x8_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4577, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4578, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4579, x0, x1, x2, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4580, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4581, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4582, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88, x89_c, x90, x91, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4583, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x52, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4584, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4585, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4586, x1, x2_c, x6, x7_c, x8, x9, x10, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4587, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x91_c, x92_c, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4588, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4589, x0_c, x3, x15_c, x16_c, x18_c, x23, x27, x33_c, x34_c, x38, x42, x43_c, x46_c, x47_c, x48_c, x51, x60, x61_c, x63, x64, x68_c, x70_c, x74_c, x79_c, x82_c, x84_c, x85_c, x86, x87, x88_c, x89_c, x90_c, x91, x99);
and (w4590, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4591, x49, x68_c, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4592, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4593, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4594, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4595, x15_c, x19, x23_c, x35, x45, x46, x60_c, x63, x69_c, x72, x79, x84, x90_c, x93);
and (w4596, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4597, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35_c, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4598, x12_c, x40, x72, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4599, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x96, x98, x99_c);
and (w4600, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4601, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4602, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x55_c, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4603, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x68, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4604, x0_c, x2_c, x6_c, x7, x8, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4605, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96, x97_c);
and (w4606, x22_c, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4607, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x73, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4608, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4609, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x92_c, x93_c, x94_c, x95, x97_c);
and (w4610, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x49, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4611, x0, x2, x3, x5, x7_c, x8, x10_c, x12_c, x13_c, x15, x17_c, x18, x19, x20, x22, x23_c, x24, x25, x26, x27_c, x28, x29, x31_c, x32_c, x35, x36, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x48_c, x49_c, x51_c, x52, x53_c, x54, x55, x56, x58, x59, x60_c, x62, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80_c, x81, x82_c, x83, x84, x85, x86, x87, x88_c, x89_c, x90, x91, x92, x93, x94, x95_c, x97, x98_c, x99);
and (w4612, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91_c, x92, x95_c, x96, x98, x99);
and (w4613, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x60_c, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4614, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x96_c, x98, x99);
and (w4615, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4616, x2_c, x10_c, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4617, x0, x1_c, x3, x4, x5, x6_c, x8_c, x9_c, x10, x12, x13_c, x14_c, x15_c, x16, x17_c, x18_c, x20, x21_c, x22, x24_c, x25, x26, x27, x28_c, x29, x30, x32, x33_c, x34_c, x36_c, x37, x39_c, x40, x41, x42, x43, x44, x45, x46, x47, x49_c, x50_c, x52_c, x55, x57_c, x58, x59_c, x60, x62_c, x63, x64, x65, x68_c, x70, x71, x72_c, x73, x75, x76_c, x78, x79_c, x80, x82_c, x83, x86, x87_c, x88, x89_c, x90, x91, x93_c, x94, x95, x97, x99_c);
and (w4618, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x47, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4619, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x67, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4620, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4621, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88_c);
and (w4622, x5, x10, x16, x21_c, x25, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w4623, x12_c, x32, x91, x99_c);
and (w4624, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71, x83_c);
and (w4625, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x70_c, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4626, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4627, x12_c, x32, x83_c, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4628, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4629, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4630, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x65, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4631, x12_c, x32, x51, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4632, x2_c, x3, x4_c, x5_c, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4633, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x73, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4634, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4635, x1, x3_c, x11_c, x13_c, x19, x20, x25, x26_c, x27, x32_c, x34_c, x41_c, x43_c, x44_c, x45, x53, x57, x59, x61, x70, x83, x88, x94, x96, x97_c);
and (w4636, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4637, x0_c, x1, x2, x3_c, x4, x5_c, x6, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4638, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51_c, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4639, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4640, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4641, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x92_c, x95, x97_c);
and (w4642, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4643, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x64, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4644, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x47_c, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4645, x0, x1_c, x3_c, x4, x5, x6_c, x7, x8_c, x9_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19, x20_c, x21, x22, x23, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32_c, x33, x34, x35_c, x37, x38, x39, x40_c, x41_c, x42_c, x43_c, x45_c, x46, x47, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x57_c, x58_c, x59, x60, x61, x62_c, x63, x64_c, x65, x66_c, x68_c, x69, x70_c, x71, x72, x73, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81_c, x83_c, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99_c);
and (w4646, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4647, x2_c, x3, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4648, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4649, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4650, x0_c, x2_c, x4_c, x7_c, x11, x12, x16, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4651, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4652, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12_c, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4653, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14_c, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4654, x11_c, x62, x69_c, x75, x92, x99);
and (w4655, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x75_c, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4656, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4657, x1, x4, x5_c, x6_c, x8_c, x11, x12, x13, x14_c, x15_c, x16, x18, x19, x20, x21_c, x23, x24_c, x25_c, x27, x28_c, x29, x30_c, x35_c, x37_c, x40_c, x41, x42_c, x46_c, x48, x49, x51_c, x52_c, x53, x54, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72, x73_c, x74, x76, x77, x78_c, x79, x80_c, x82_c, x83, x84, x85, x86_c, x87_c, x91_c, x92_c, x93, x94, x96, x97_c, x98_c, x99);
and (w4658, x1, x2, x5, x6_c, x7_c, x8, x9_c, x10_c, x11, x12, x13_c, x14, x16_c, x18, x20, x21, x22_c, x24_c, x26, x27, x30_c, x31, x32, x33, x35, x37_c, x38_c, x40_c, x42, x43_c, x46_c, x47, x48_c, x49_c, x52_c, x55_c, x57, x59, x60_c, x61_c, x62_c, x63, x64_c, x66, x67, x68_c, x69, x72_c, x73, x75_c, x78, x79, x80, x82_c, x83_c, x84, x86, x87_c, x91, x93, x94, x95, x96_c, x97, x98_c, x99);
and (w4659, x0, x4, x5, x7, x9_c, x10, x14, x16, x17, x23, x24_c, x25_c, x32_c, x33_c, x40, x41, x46_c, x48, x51, x55_c, x58, x63_c, x70, x75, x79, x80_c, x85_c, x87_c, x88, x91, x94, x96);
and (w4660, x0, x3, x5, x6, x9, x10, x11_c, x14, x15_c, x18_c, x20, x21, x25_c, x26_c, x27_c, x28_c, x29, x31, x37_c, x38_c, x39_c, x42_c, x43, x44_c, x50, x51_c, x52, x53_c, x57, x58, x62_c, x63, x64, x67_c, x69, x71_c, x73_c, x74, x75_c, x81_c, x82, x83_c, x86_c, x87, x88_c, x89, x90, x92_c, x96_c, x97_c);
and (w4661, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x76, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4662, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4663, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4664, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4665, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4666, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x74_c, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w4667, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47, x82, x90_c, x96, x98, x99_c);
and (w4668, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4669, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x56_c, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4670, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4671, x12_c, x40, x45_c, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4672, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4673, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4674, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4675, x0, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4676, x5_c, x9, x27, x61_c, x76, x88_c, x91_c, x92, x95, x97_c);
and (w4677, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x53_c, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4678, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x35_c, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4679, x1, x3, x4, x5, x10_c, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4680, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91, x92, x93_c, x94_c, x95, x97_c, x98, x99_c);
and (w4681, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
assign w4682 = x34;
and (w4683, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x55_c, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4684, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4685, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4686, x0, x1, x2_c, x4_c, x7_c, x10_c, x13_c, x15_c, x18_c, x20_c, x23_c, x27_c, x28, x29_c, x31, x35, x37, x41, x42, x44_c, x46, x48_c, x49_c, x50, x55_c, x56_c, x57, x58_c, x60_c, x64, x66, x68_c, x73_c, x74, x75_c, x76_c, x78, x79_c, x82, x83, x85_c, x86_c, x90_c, x93, x94, x95_c);
and (w4687, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c, x98_c, x99);
and (w4688, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x79, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4689, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x39, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4690, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4691, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4692, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4693, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x91_c, x93_c, x94_c, x95_c, x97, x98, x99_c);
and (w4694, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x66_c, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4695, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x80, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4696, x8, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4697, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7, x8, x9_c, x10_c, x11, x12, x13_c, x14_c, x15, x16_c, x17_c, x18, x20_c, x21_c, x22_c, x23_c, x25_c, x26, x27_c, x28, x29, x30_c, x31_c, x32, x33, x34_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x41, x42, x43_c, x44_c, x45, x46_c, x47_c, x48, x49, x51, x52, x53, x54_c, x55, x56_c, x57_c, x58, x59_c, x60_c, x61_c, x62, x64_c, x65_c, x66_c, x67_c, x68, x69, x70, x71_c, x72, x73_c, x74, x75, x76_c, x77, x78_c, x79_c, x80_c, x81_c, x82, x83, x84, x85, x86_c, x87, x88, x89, x90_c, x91, x92_c, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w4698, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4699, x0_c, x5, x23_c, x30_c, x31, x32_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4700, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4701, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x78_c, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4702, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4703, x1_c, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4704, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4705, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x77_c, x82, x83, x93_c, x97_c);
and (w4706, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4707, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4708, x2_c, x11, x20, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4709, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77_c, x81_c, x82, x88_c, x93_c, x95_c);
and (w4710, x1_c, x2, x4, x5, x6_c, x9_c, x10, x11, x12_c, x14_c, x17, x18_c, x20_c, x21, x22_c, x25, x26_c, x28, x30, x31_c, x32, x34_c, x35_c, x37, x38, x42_c, x46, x47, x48_c, x52_c, x54_c, x57, x59_c, x60, x64_c, x66, x67, x68, x70_c, x73, x75_c, x77, x84_c, x85, x86, x87_c, x88, x90_c, x91, x94, x95_c, x98_c, x99_c);
and (w4711, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x12_c, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4712, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4713, x13_c, x14_c, x37_c, x39_c, x45_c, x53, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4714, x0, x13_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4715, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79, x81, x84, x85, x95, x99);
and (w4716, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x33, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4717, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92_c, x93_c, x97_c);
and (w4718, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4719, x12_c, x29, x46, x47_c, x48_c, x50_c, x61_c, x66, x67_c, x77, x78, x94);
and (w4720, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x89_c, x91_c, x92, x93, x94, x95, x96, x97_c, x99_c);
and (w4721, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x16, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4722, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4723, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4724, x0_c, x1_c, x2_c, x3, x5, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14, x15, x17_c, x18, x20, x21, x22_c, x23_c, x24_c, x25, x28, x29, x31, x32_c, x33_c, x34, x35, x36, x37, x38, x39, x40, x41, x42_c, x43_c, x44_c, x45, x46_c, x47, x48_c, x49, x50_c, x51, x53, x54, x56, x58_c, x60_c, x61_c, x62_c, x63_c, x65_c, x66_c, x68, x69_c, x70_c, x71_c, x73_c, x74_c, x75, x76_c, x77_c, x78_c, x79, x82, x83_c, x84, x86, x87, x88, x89_c, x91, x93, x94_c, x95, x96_c, x97_c, x98, x99);
and (w4725, x2_c, x3, x4, x6_c, x11, x12, x13, x15, x16_c, x20_c, x22, x23, x24_c, x25, x32_c, x33_c, x34_c, x38, x39_c, x43_c, x45, x46_c, x49_c, x50, x56, x57_c, x58, x59, x62_c, x64_c, x66, x67_c, x70_c, x73, x74_c, x79, x80, x83_c, x84, x85_c, x86, x90_c, x91, x93_c, x94);
and (w4726, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x52, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4727, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4728, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x92, x96_c, x97);
and (w4729, x8, x21_c, x25_c, x27_c, x33_c, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4730, x0, x1, x2_c, x3_c, x5_c, x9, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4731, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4732, x12_c, x32, x45_c, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4733, x0, x7_c, x9, x12, x21_c, x34, x36_c, x39_c, x44_c, x49, x50, x52_c, x60_c, x66, x75, x76_c, x80, x81_c, x82_c, x86, x92_c, x93);
and (w4734, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x23, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4735, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4736, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x37, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4737, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4738, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4739, x6, x17_c, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4740, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4741, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4742, x0_c, x5_c, x15, x18, x19, x22, x31, x36, x39_c, x41, x47_c, x49_c, x51, x61, x64, x67, x77, x80_c, x88, x91_c, x96);
and (w4743, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96_c, x97_c);
and (w4744, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w4745, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93, x95, x97_c);
and (w4746, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x71, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4747, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4748, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x20, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w4749, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4750, x0, x6_c, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w4751, x0, x1, x2_c, x3, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4752, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x62, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4753, x3, x7_c, x8_c, x13_c, x17_c, x19, x21_c, x26, x29, x38_c, x39, x42, x45, x47, x57, x62, x75_c, x80_c, x81, x86, x90, x93, x94, x96_c, x97, x99_c);
and (w4754, x49, x50_c, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4755, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4756, x28_c, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4757, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4758, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4759, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4760, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x20_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4761, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x83_c, x93_c, x97_c);
and (w4762, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97, x98, x99);
and (w4763, x9, x12, x13_c, x14_c, x23_c, x31_c, x32_c, x43_c, x45_c, x48, x51_c, x52_c, x54, x55, x68, x87_c, x94, x95, x96_c);
and (w4764, x0_c, x3_c, x10, x15, x16_c, x19_c, x20_c, x22_c, x23, x27, x29, x30, x33, x34, x35, x42, x43_c, x53_c, x57_c, x60_c, x62_c, x63, x64_c, x69, x71_c, x72_c, x75, x77, x79, x80, x85, x86_c, x93, x96_c);
and (w4765, x3_c, x6_c, x8_c, x11_c, x12_c, x16_c, x18, x21, x23, x25_c, x32, x33, x34_c, x36, x43_c, x46, x52, x53, x58, x59_c, x60, x62_c, x64, x66_c, x71_c, x72_c, x79, x80, x81_c, x88_c, x90_c, x92, x98_c);
and (w4766, x1, x2_c, x5, x7_c, x8, x9_c, x10_c, x12_c, x13, x16, x17_c, x18_c, x19, x20_c, x21, x22_c, x23_c, x24_c, x25, x26_c, x27_c, x28_c, x30_c, x31_c, x32_c, x38_c, x40_c, x41, x42_c, x44_c, x45_c, x48, x51_c, x52_c, x53_c, x54, x55, x56, x61, x62_c, x63_c, x64, x65, x66, x68, x69, x72, x73, x74, x75_c, x78, x80_c, x81, x82_c, x84, x85_c, x87, x88, x89, x90_c, x91, x92_c, x93, x97, x99);
and (w4767, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4768, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4769, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91_c, x93_c, x97_c);
and (w4770, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92, x95, x96, x97_c, x98, x99_c);
and (w4771, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4772, x0, x1_c, x2, x3, x4_c, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x13_c, x14, x15_c, x17, x18_c, x19_c, x20, x21_c, x22, x23, x24, x25, x26, x27, x28, x29_c, x30_c, x31, x32, x33, x34_c, x35, x36, x37_c, x39, x40_c, x41, x42_c, x43, x44, x45_c, x46_c, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57_c, x58, x59, x60, x61, x62, x63_c, x64, x65, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x72, x73, x74_c, x75, x76_c, x77, x78, x79, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87_c, x88_c, x89_c, x90, x91_c, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98_c, x99);
and (w4773, x3, x13, x24, x27_c, x29, x31_c, x33_c, x34_c, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4774, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82_c, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4775, x12_c, x32, x82, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4776, x2_c, x52_c, x70_c);
and (w4777, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4778, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x68_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4779, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60_c, x82, x90_c, x96, x98, x99_c);
and (w4780, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x68_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4781, x2_c, x4, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4782, x0, x1_c, x2, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4783, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4784, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98_c, x99_c);
and (w4785, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x66, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4786, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4787, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x88_c, x89, x90, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4788, x0_c, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4789, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71_c, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4790, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4791, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74_c, x76, x85, x89, x93, x97_c);
and (w4792, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88, x90_c, x92, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4793, x2_c, x11, x29_c, x95, x96, x98, x99);
and (w4794, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x30, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4795, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4796, x5, x10, x16, x21_c, x34_c, x35, x41, x42, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w4797, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x69, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4798, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4799, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x54_c, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4800, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x75_c, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4801, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4802, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c, x99);
and (w4803, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4804, x13_c, x14_c, x37_c, x39_c, x41_c, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4805, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4806, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67_c, x83_c);
and (w4807, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w4808, x12_c, x40, x69, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4809, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96_c);
and (w4810, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4811, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x30, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4812, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86_c, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4813, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41_c, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4814, x2_c, x4, x6, x7_c, x10_c, x11_c, x13, x17, x18, x30_c, x31, x38, x40_c, x41, x43, x48, x50, x52, x53_c, x55, x57, x63, x65_c, x68, x69, x72, x75, x77, x79, x84_c, x85, x89, x92, x94_c, x95_c, x97, x99_c);
and (w4815, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4816, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4817, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36_c, x40, x82, x90_c, x96, x98, x99_c);
and (w4818, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4819, x5_c, x9, x13, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4820, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4821, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4822, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4823, x4_c, x5, x83_c);
and (w4824, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x71_c, x81_c, x82, x88_c, x93_c, x95_c);
and (w4825, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x39_c, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4826, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81, x83_c);
and (w4827, x12_c, x32, x37, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4828, x0_c, x2_c, x3, x4, x5, x7, x9, x10_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4829, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x18, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4830, x10_c, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w4831, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x88, x90_c, x91, x92, x95, x97_c);
and (w4832, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91_c, x92_c, x93_c, x95_c, x96, x98, x99);
and (w4833, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4834, x0_c, x2_c, x3, x5_c, x6, x7, x9, x10_c, x11, x13, x14_c, x15, x16, x17, x18, x19, x21, x22, x25_c, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x35, x37_c, x39_c, x40, x42_c, x43, x44, x45_c, x47, x48_c, x49_c, x50_c, x51, x53, x54_c, x55_c, x56_c, x57, x58, x60, x61, x62_c, x63_c, x64_c, x65_c, x67_c, x68, x69, x70, x71_c, x72, x73_c, x75_c, x76, x77_c, x79_c, x81, x83, x84, x85_c, x87_c, x88, x90, x92_c, x93_c, x94, x95, x96_c, x99_c);
and (w4835, x0, x1, x2, x3_c, x5_c, x8_c, x9, x10_c, x14, x16, x17, x18, x21_c, x22, x24, x25_c, x26, x30_c, x31, x32, x33, x34_c, x36, x38_c, x39_c, x40, x41_c, x42_c, x45, x46, x47, x48_c, x49, x50, x51, x53, x54, x55, x57, x60, x61, x62, x64_c, x66_c, x69, x70_c, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80, x81, x82_c, x83, x90, x91, x92, x93_c, x94, x96_c, x97, x99);
and (w4836, x12_c, x40, x82, x83_c, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4837, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4838, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4839, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x95, x96_c, x97_c, x98, x99_c);
and (w4840, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x29_c, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4841, x0, x1, x2, x3_c, x4, x5, x6, x7_c, x8_c, x9, x10, x12, x13, x14, x15, x17_c, x18, x19, x20_c, x21, x24_c, x25_c, x26_c, x27_c, x32, x33_c, x34_c, x35, x36, x38, x40_c, x42_c, x45_c, x46, x47, x49_c, x50_c, x51_c, x54_c, x59_c, x60, x61, x63, x64, x65, x66_c, x68_c, x70_c, x71_c, x72_c, x73_c, x74, x76, x77_c, x78, x79_c, x80, x83, x87_c, x88_c, x89_c, x90, x92, x94_c, x97_c, x99_c);
and (w4842, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4843, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x69_c, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4844, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4845, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4846, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43_c, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4847, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4848, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4849, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4850, x12_c, x40, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4851, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x40, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4852, x3_c, x6_c, x7_c, x15_c, x21, x27_c, x29_c, x32_c, x34, x36, x37, x41, x42, x48_c, x57_c, x66_c, x68, x76, x77_c, x78_c, x83_c, x93_c, x98);
and (w4853, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x56_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4854, x12_c, x32, x81, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4855, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4856, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4857, x13_c, x24, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w4858, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x39_c, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4859, x0_c, x1_c, x2_c, x3, x4, x5, x6_c, x7_c, x8, x9_c, x10, x11, x13, x14, x16, x17_c, x20, x21, x23, x24, x27, x28, x29, x32, x34, x35_c, x36_c, x37, x38_c, x39_c, x42, x43, x46_c, x47, x48_c, x49, x50, x51_c, x52, x53_c, x54, x55, x56_c, x58, x59, x60, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69_c, x70, x72_c, x76, x78_c, x79_c, x80, x82, x83_c, x85_c, x87, x89, x90_c, x91_c, x92_c, x93, x94_c, x95, x96, x98, x99);
and (w4860, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w4861, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4862, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x35, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4863, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x84_c, x85_c, x97_c, x98_c, x99_c);
and (w4864, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x70, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4865, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x90_c, x92_c, x94, x96_c, x97, x99);
and (w4866, x0, x1, x2, x3_c, x4, x5, x6, x7_c, x9_c, x10_c, x11, x12, x14, x17_c, x18_c, x19_c, x20_c, x21_c, x22, x23_c, x24, x25_c, x28_c, x29, x31_c, x35, x36, x37_c, x38_c, x39, x42, x43, x44, x46_c, x47, x48_c, x49_c, x50_c, x51, x52_c, x53_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x70_c, x72_c, x74, x75, x77, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x85_c, x86, x88_c, x89, x90, x92_c, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w4867, x1, x12_c, x21, x51, x64, x74_c, x78_c, x96_c);
and (w4868, x5, x10, x16, x21_c, x23, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4869, x6_c, x7, x8_c, x12_c, x13, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4870, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4871, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4872, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4873, x0_c, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x11, x12_c, x13, x14_c, x15_c, x16, x17, x18, x19_c, x20_c, x22_c, x23_c, x24_c, x25_c, x26_c, x28, x29_c, x30, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37, x38_c, x39, x40, x41_c, x42_c, x43, x44, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x54, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63, x64_c, x65, x68_c, x69, x70_c, x73, x74, x75, x76, x77, x78_c, x79_c, x80, x81_c, x82, x83, x85_c, x86, x87, x88, x89_c, x90_c, x91, x92_c, x94, x95, x96_c, x97, x98, x99);
and (w4874, x0_c, x5, x23_c, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4875, x12_c, x32, x91, x98_c, x99);
and (w4876, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x32_c, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4877, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x61, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w4878, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4879, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4880, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4881, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x75, x77, x82, x83, x93_c, x97_c);
and (w4882, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4883, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59, x83_c);
and (w4884, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x84_c, x85_c, x97_c, x99);
and (w4885, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4886, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4887, x0_c, x1, x2, x3, x4, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12, x13, x14, x15_c, x16_c, x17_c, x18, x19, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x32, x34_c, x35, x36, x38_c, x39, x40_c, x41_c, x42, x43_c, x44, x45, x46_c, x47, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x57_c, x58_c, x59, x60_c, x61, x62, x63_c, x64_c, x65_c, x66, x67, x68, x69, x70, x71_c, x72, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92, x93, x94, x96, x98, x99);
and (w4888, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x28, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4889, x0, x1_c, x3_c, x7_c, x8_c, x9_c, x10, x11, x12, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x30_c, x31_c, x32, x33, x34, x35_c, x36, x37, x38_c, x39_c, x40, x41_c, x42_c, x43, x45, x47_c, x48, x49_c, x50, x51, x52, x53_c, x54_c, x55, x56_c, x57_c, x58_c, x59, x61_c, x63, x64, x65_c, x66, x67_c, x68, x69, x70, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78_c, x79, x80_c, x81, x82_c, x83_c, x84, x85, x86, x88, x89, x90, x91, x92_c, x93_c, x94, x95, x96_c, x97, x98);
and (w4890, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4891, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17_c, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4892, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91_c, x93_c, x95_c, x96, x98, x99);
and (w4893, x4_c, x10, x15_c, x22_c, x24_c, x25, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4894, x9, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4895, x26_c, x28_c, x40_c, x44, x57_c, x62, x71_c);
and (w4896, x7, x12, x14_c, x18, x20, x28_c, x35_c, x36_c, x38, x43, x55_c, x63_c, x74_c, x80, x85_c, x87, x89_c, x91, x92, x94, x95);
and (w4897, x2_c, x3, x4, x7, x11_c, x13_c, x16, x18_c, x19_c, x21_c, x26, x35, x37, x38_c, x41, x44_c, x52_c, x56, x57, x60_c, x62, x68, x70, x75_c, x76, x82_c, x83, x91, x96, x98);
and (w4898, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x57, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4899, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4900, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x22, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4901, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4902, x0_c, x2, x3_c, x4, x5, x6, x7_c, x9_c, x10_c, x13, x14, x15, x17_c, x18, x19, x21_c, x23, x24, x25_c, x26_c, x27, x29_c, x30, x32, x33_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41, x42, x43, x44_c, x45, x46, x47, x48_c, x50, x51, x52, x53_c, x54_c, x55, x58, x59_c, x60_c, x61_c, x62, x63, x64, x65_c, x66_c, x67_c, x68_c, x70_c, x71_c, x73_c, x74_c, x75_c, x77_c, x78, x79, x80_c, x81_c, x82, x83_c, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91, x94, x95, x97_c, x98, x99);
and (w4903, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w4904, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w4905, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x68_c, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w4906, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x42, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4907, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x88_c, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4908, x2_c, x4, x5_c, x9, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4909, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4910, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4911, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4912, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4913, x0_c, x5, x23, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4914, x0, x1_c, x3, x4_c, x6_c, x8_c, x12_c, x14, x20_c, x23, x24_c, x26_c, x29_c, x31_c, x32_c, x34, x36, x38, x40, x41_c, x43, x47, x52_c, x55_c, x58, x64_c, x66, x70, x74_c, x78_c, x79_c, x81, x84_c, x86_c, x92, x94, x98_c, x99);
and (w4915, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x96, x98, x99);
and (w4916, x0_c, x1, x5, x7_c, x8, x9_c, x10, x11, x12, x13, x14_c, x16_c, x17, x19, x21_c, x22_c, x23, x24, x26, x27_c, x28, x30, x31, x32_c, x34, x35, x36, x37, x38, x39_c, x40, x41, x42, x44_c, x46, x47_c, x48, x49, x50_c, x51, x52_c, x53_c, x54_c, x55, x56, x57, x58, x59, x60, x61_c, x62, x63, x64, x65_c, x67, x68, x69, x71_c, x72_c, x74_c, x78_c, x79_c, x80_c, x81, x82_c, x83_c, x84, x85, x86, x87_c, x88, x89_c, x90_c, x91, x92, x95_c, x96_c, x97_c, x99_c);
and (w4917, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x87_c, x89, x93_c, x95_c, x96_c, x97_c);
and (w4918, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4919, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x26, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4920, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x21_c, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4921, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w4922, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w4923, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x74, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4924, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4925, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87, x90_c, x93_c, x97_c);
and (w4926, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4927, x3_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w4928, x0, x6, x7_c, x9, x10, x15_c, x32_c, x36, x51_c, x63, x69_c, x70, x72, x78_c, x89_c, x92_c, x97);
and (w4929, x12_c, x32, x49_c, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w4930, x0, x2, x3, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4931, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4932, x5_c, x7, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4933, x0_c, x2_c, x3_c, x4, x6, x7, x8, x11_c, x13, x14, x15_c, x16, x17, x18, x21_c, x26_c, x27, x28, x30_c, x31_c, x32, x34, x35, x36_c, x38, x40, x43, x47_c, x48_c, x53, x54, x55_c, x57, x58_c, x63_c, x65_c, x66, x68_c, x69, x70_c, x71, x75, x76, x77, x78_c, x79, x80_c, x83_c, x84_c, x85, x87_c, x90, x92, x93_c, x97_c, x98, x99_c);
and (w4934, x0_c, x5, x21, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4935, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x91_c, x92, x95, x97_c);
and (w4936, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x43_c, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4937, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4938, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4939, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4940, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4941, x2, x4_c, x5, x6, x7_c, x9_c, x12_c, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4942, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4943, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w4944, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4945, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4946, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77_c, x81, x84, x85, x95, x99);
and (w4947, x12_c, x40, x59_c, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4948, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32_c, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4949, x0_c, x1, x2, x3_c, x4_c, x5, x6_c, x7_c, x8, x9_c, x11_c, x13, x14_c, x15, x17, x18, x19_c, x25_c, x26_c, x27_c, x28_c, x29_c, x30, x31_c, x32_c, x33_c, x35, x37_c, x38_c, x39, x40, x41, x42, x43_c, x44_c, x45, x47_c, x48, x49_c, x51_c, x52, x53_c, x54_c, x56_c, x57, x58_c, x59_c, x60_c, x61, x63_c, x64, x67, x68, x69, x70, x71_c, x72_c, x73_c, x74, x75, x77_c, x78_c, x79_c, x80_c, x81_c, x83, x84, x87_c, x88, x89_c, x90, x91_c, x92, x95, x96, x99);
and (w4950, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4951, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4952, x3, x6, x8_c, x10, x12_c, x14_c, x16, x19_c, x25, x34, x35_c, x38_c, x39_c, x40_c, x41, x42, x45_c, x46_c, x47_c, x48, x51, x53_c, x56_c, x59, x60_c, x63_c, x65_c, x70, x73, x75, x76, x77, x78, x79, x81, x83_c, x86_c, x89_c, x95_c, x97_c);
and (w4953, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w4954, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x79, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4955, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4956, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4957, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x20, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w4958, x9_c, x17_c, x26, x27, x28_c, x32, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4959, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4960, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4961, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4962, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4963, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x22, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4964, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w4965, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4966, x12_c, x40, x79, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w4967, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w4968, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4969, x0, x1, x2, x5, x6, x7_c, x9_c, x10_c, x11_c, x12, x13, x14_c, x16_c, x17_c, x20_c, x21, x24, x25, x26, x27, x29, x31_c, x32_c, x33, x34_c, x37, x38, x40, x41_c, x42_c, x43, x44_c, x46_c, x48, x49, x50, x51_c, x53, x54, x55_c, x57_c, x58, x60, x61_c, x62_c, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x74_c, x75, x76, x77_c, x78_c, x79, x80_c, x81, x82_c, x86_c, x87_c, x88, x89, x90, x91_c, x92, x93, x94, x95, x97_c, x98);
and (w4970, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w4971, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x30, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4972, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w4973, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x90_c, x91, x96, x97, x99);
and (w4974, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w4975, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x55_c, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w4976, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x16_c, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4977, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x29_c, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4978, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x74_c, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w4979, x73, x95, x96, x98, x99);
and (w4980, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x89_c, x91, x93, x97_c);
and (w4981, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4982, x8, x21_c, x25_c, x27_c, x28, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4983, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x68, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4984, x13_c, x49, x64, x71, x72_c, x75_c, x81_c, x87, x90, x93_c, x97_c);
and (w4985, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4986, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19_c, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w4987, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x56_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w4988, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x94, x95, x96_c, x97, x98, x99_c);
and (w4989, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4990, x0_c, x5, x21, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4991, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4992, x0_c, x1_c, x3, x4, x5, x7, x8_c, x10_c, x13, x16_c, x18, x19, x20, x22, x24, x25_c, x26_c, x28_c, x29_c, x30, x33_c, x35, x36, x38, x39, x40, x41_c, x43, x44_c, x45_c, x46_c, x50_c, x52, x53_c, x54_c, x57, x58_c, x60_c, x61_c, x62, x64_c, x65, x68_c, x70, x71_c, x72, x73_c, x74, x75_c, x76, x81_c, x83_c, x85, x86, x87_c, x89, x94, x95_c, x96_c);
and (w4993, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90, x93_c, x95_c);
and (w4994, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79, x85, x89, x93, x97_c);
and (w4995, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89_c);
and (w4996, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w4997, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w4998, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w4999, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5000, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x53_c, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5001, x5_c, x9, x27, x49, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5002, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5003, x0, x1, x2, x4, x6, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5004, x12_c, x32, x73, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5005, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5006, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5007, x5, x8_c, x10_c, x11, x14, x21, x22_c, x28, x32_c, x33, x47, x49_c, x51, x57, x63, x67_c, x74_c, x77, x80_c, x84, x88, x94);
and (w5008, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x90_c, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5009, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5010, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94, x95_c, x96, x98, x99);
and (w5011, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x93, x95_c, x96, x98, x99);
and (w5012, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w5013, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97, x98, x99);
and (w5014, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x97_c, x98, x99_c);
and (w5015, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x97_c);
and (w5016, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5017, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5018, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79, x82, x83, x93_c, x97_c);
and (w5019, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x77_c, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5020, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5021, x0_c, x1_c, x3, x4_c, x5, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5022, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5023, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45_c, x82, x90_c, x96, x98, x99_c);
and (w5024, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5025, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5026, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91_c, x93_c, x97_c);
and (w5027, x0, x1, x2_c, x3, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5028, x0_c, x2_c, x21_c, x34_c, x38, x60, x78, x83, x84, x86_c, x87);
and (w5029, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5030, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x93_c, x97, x98, x99_c);
and (w5031, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45, x83_c);
and (w5032, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x12_c, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5033, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x75, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5034, x4, x5, x7_c, x10_c, x11_c, x18, x19, x21_c, x22, x28, x29, x30, x31_c, x32_c, x35_c, x36, x37_c, x38, x45_c, x49, x51, x52, x53_c, x55, x59, x62_c, x64_c, x67, x69_c, x70, x74_c, x75, x78, x79, x80_c, x81, x83_c, x86_c, x87_c, x90, x94, x95, x96, x97);
and (w5035, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5036, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5037, x0, x1, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5038, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5039, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x69, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5040, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5041, x4, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w5042, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x45_c, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5043, x13_c, x49, x64_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w5044, x12, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5045, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x41_c, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w5046, x5_c, x6, x7, x8, x9_c, x12_c, x14, x16_c, x17_c, x18, x19, x22_c, x23_c, x26, x30, x31_c, x33, x34, x36, x40, x47_c, x48, x53, x54_c, x57_c, x58, x61_c, x62, x65_c, x66, x68_c, x69_c, x70, x71, x72, x73_c, x75_c, x81_c, x86_c, x88, x89_c, x91, x92_c, x93_c, x98_c);
and (w5047, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x50_c, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5048, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44, x82, x90_c, x96, x98, x99_c);
and (w5049, x2, x4_c, x6_c, x7_c, x12_c, x13, x20, x23_c, x35, x36_c, x47, x50, x51, x70_c, x78_c, x90_c, x96);
and (w5050, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5051, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5052, x0_c, x1, x2_c, x3_c, x4_c, x5, x6_c, x7_c, x8, x9, x10_c, x12, x13_c, x15_c, x17_c, x19, x20, x21_c, x22, x23_c, x24, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34, x35, x36_c, x37, x38, x39_c, x40, x42_c, x43_c, x44_c, x45_c, x46, x47, x48_c, x49_c, x50, x51_c, x52, x53, x54, x55, x56_c, x57, x58, x59, x61, x62_c, x63_c, x64, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x83, x84, x85_c, x86_c, x87, x88, x89_c, x90_c, x91_c, x92_c, x94_c, x95_c, x96, x97_c, x98, x99_c);
and (w5053, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5054, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5055, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13_c, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5056, x0, x2, x3, x4, x7, x10, x13_c, x14_c, x17_c, x19, x20, x21, x24, x25, x27_c, x28_c, x29, x30_c, x31_c, x32_c, x33_c, x35_c, x36_c, x40, x41, x42_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x52_c, x54, x56, x57_c, x58, x59_c, x60_c, x62_c, x64_c, x65_c, x66, x67, x69_c, x70_c, x72_c, x73, x74, x75, x77_c, x78_c, x79_c, x80, x81, x82, x83_c, x84_c, x85_c, x86, x87_c, x88_c, x89_c, x91_c, x92, x93_c, x94, x95_c, x96, x97_c, x98, x99);
and (w5057, x53_c, x83_c);
and (w5058, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98_c);
and (w5059, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78_c, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5060, x12_c, x40, x82, x89, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5061, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5062, x0_c, x3_c, x6, x7, x8_c, x9_c, x12_c, x13_c, x14_c, x15, x16, x19, x20_c, x21_c, x22_c, x24, x25, x26_c, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x38_c, x39, x41, x42_c, x43, x45, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x54, x55_c, x57_c, x58_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x67, x68_c, x70, x71_c, x72, x75, x76, x77_c, x78, x79_c, x80_c, x85_c, x87, x89, x91_c, x92, x93, x94, x95_c, x96, x97, x98, x99);
and (w5063, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5064, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5065, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x37_c, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5066, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54_c, x82, x90_c, x96, x98, x99_c);
and (w5067, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5068, x4_c, x7_c, x13, x18_c, x19_c, x20, x21_c, x23_c, x25, x30_c, x32_c, x37_c, x59, x67, x68_c, x73_c, x74_c, x88_c, x93, x94_c, x95);
and (w5069, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x95_c, x96_c, x97);
and (w5070, x2_c, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5071, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5072, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42_c, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5073, x0, x3_c, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5074, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x93_c, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w5075, x1, x7, x8_c, x10, x17_c, x23, x26_c, x34, x40, x46, x48_c, x49_c, x58_c, x61_c, x62, x68_c, x69, x72, x74, x80_c);
and (w5076, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5077, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8, x9, x13, x14, x15_c, x17_c, x18_c, x19, x21, x22_c, x23_c, x24, x25_c, x26, x27_c, x28_c, x29_c, x31_c, x33_c, x35, x36_c, x38, x39_c, x40_c, x42_c, x43, x46_c, x47, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56, x57, x58, x59_c, x60_c, x61_c, x63_c, x64, x66, x67, x68, x69_c, x70, x71_c, x72_c, x73_c, x74, x75, x77_c, x78_c, x83, x85_c, x86, x88, x90, x91_c, x93_c, x95, x96, x97_c, x98, x99_c);
and (w5078, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x38_c, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5079, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97, x99);
and (w5080, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5081, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5082, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5083, x1_c, x2, x4_c, x6_c, x10, x13_c, x14_c, x19_c, x20, x21_c, x23, x24_c, x28_c, x29, x31, x34_c, x35_c, x36_c, x40_c, x42, x47_c, x48_c, x49, x50, x51_c, x53_c, x54, x55, x57_c, x58_c, x61_c, x62_c, x63_c, x65, x66_c, x67, x69_c, x70, x71, x73, x75, x76_c, x77, x80, x82_c, x83_c, x84, x85_c, x86, x89, x95);
and (w5084, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x47, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5085, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5086, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5087, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x29, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5088, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5089, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5090, x1, x4_c, x5_c, x6, x7_c, x8_c, x11, x12_c, x13_c, x15, x16, x20, x22, x26_c, x28, x30_c, x32_c, x34_c, x35_c, x36, x37_c, x43_c, x44, x45, x47_c, x49_c, x51, x53, x54_c, x56_c, x57, x58, x59_c, x60, x61, x62_c, x66_c, x67, x68, x72_c, x73_c, x78, x83, x84_c, x85, x86_c, x87_c, x88_c, x89_c, x92_c, x93_c, x96, x97, x99);
and (w5091, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x45, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5092, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5093, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5094, x1, x3_c, x4_c, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12, x13_c, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x28_c, x29_c, x30, x31, x32, x33, x39, x40, x42_c, x44, x45_c, x46_c, x47, x48, x49, x50, x51, x52_c, x54_c, x55, x56_c, x57_c, x58_c, x60_c, x61_c, x62, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x73_c, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83, x84_c, x85, x86_c, x87, x88, x89, x90_c, x91, x92_c, x93, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w5095, x3, x5, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5096, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x68, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5097, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64, x73_c, x76, x85, x89, x93, x97_c);
and (w5098, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5099, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5100, x0_c, x2_c, x14_c, x17, x18, x28, x30_c, x33, x36, x37_c, x40, x45_c, x49_c, x50, x60, x69_c, x71, x72, x75_c, x82, x85, x97);
and (w5101, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x74, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5102, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5103, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5104, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x39_c, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5105, x1, x3_c, x7, x8_c, x9, x10_c, x12_c, x13_c, x14, x19_c, x21_c, x22_c, x24, x25, x27, x28_c, x30, x31_c, x36_c, x37_c, x38_c, x41, x42, x44, x47, x52_c, x53, x54_c, x55_c, x56, x59, x60, x65, x66_c, x73_c, x75_c, x78_c, x79_c, x81_c, x82_c, x83_c, x85, x86_c, x89_c, x90_c, x91, x99_c);
and (w5106, x0_c, x1_c, x2_c, x3, x4_c, x5, x6_c, x9, x10_c, x13_c, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x27, x28, x29, x30_c, x31_c, x33, x34, x35_c, x36, x37, x38_c, x39, x40_c, x41_c, x42_c, x44_c, x45, x46, x47, x48_c, x49_c, x53_c, x54, x55, x56, x57_c, x58, x59_c, x60, x61_c, x64_c, x67_c, x68_c, x69_c, x70_c, x72, x73, x74_c, x76, x77_c, x78, x79, x81, x82_c, x83_c, x84, x85, x86, x88_c, x89_c, x92_c, x93_c, x94, x95_c, x96_c, x99_c);
and (w5107, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5108, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5109, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5110, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79_c);
and (w5111, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x98_c, x99);
and (w5112, x27_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5113, x7, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w5114, x49, x64_c, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5115, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5116, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5117, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5118, x1, x4, x7, x8_c, x11, x12, x13, x14, x19_c, x21, x22_c, x24, x27, x28_c, x38, x43_c, x53_c, x54, x55_c, x56_c, x59_c, x69_c, x72_c, x73_c, x74, x77, x83_c, x84, x85_c, x96_c, x98_c);
and (w5119, x6_c, x7_c, x8_c, x9, x10, x14_c, x15_c, x20, x21, x22, x26_c, x27, x28, x29_c, x30, x31_c, x32_c, x35_c, x37_c, x38_c, x40_c, x41_c, x42_c, x43_c, x47_c, x48, x51, x53_c, x54, x56, x57_c, x60, x64_c, x65_c, x66, x71_c, x73, x74_c, x75, x77_c, x79_c, x80, x81, x82, x84_c, x86_c, x87_c, x88, x89_c, x92_c, x93_c, x94_c, x95_c, x96_c, x99);
and (w5120, x0_c, x3_c, x4_c, x6, x7, x8_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5121, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x56, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5122, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5123, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98);
and (w5124, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x96, x98, x99_c);
and (w5125, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5126, x1, x3_c, x6_c, x19_c, x26, x27, x29, x30, x33_c, x39_c, x40, x41, x45_c, x47_c, x52, x58_c, x62_c, x67, x70, x72, x74, x87_c, x88_c, x91_c, x94, x95_c, x97_c, x98_c);
and (w5127, x0_c, x8_c, x9, x11_c, x13_c, x14, x17, x18, x22_c, x24_c, x27_c, x30_c, x31_c, x32_c, x35_c, x37_c, x38, x54, x56_c, x58_c, x66, x67, x68, x71_c, x74_c, x77, x82_c, x84_c, x86, x87, x91_c, x98);
and (w5128, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x87, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5129, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x87, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5130, x2_c, x11, x27, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5131, x0_c, x5, x8, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5132, x0_c, x2_c, x3, x5_c, x9, x10, x11_c, x12_c, x15, x16_c, x17, x18_c, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x28_c, x30, x31, x32_c, x33_c, x35_c, x36_c, x37_c, x39_c, x42_c, x43, x45_c, x49_c, x51, x53, x57, x60_c, x61_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x71_c, x74, x76, x77_c, x79_c, x80, x82, x84_c, x85_c, x87, x93);
and (w5133, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48_c, x82, x90_c, x96, x98, x99_c);
and (w5134, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x24, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5135, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82, x85, x89, x93, x97_c);
and (w5136, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5137, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x90, x93_c, x95_c, x96, x98, x99);
and (w5138, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5139, x0, x6, x14_c, x16, x18, x19_c, x20, x22_c, x24, x25_c, x32_c, x41_c, x43_c, x46_c, x48_c, x49, x51, x55_c, x59_c, x61_c, x66, x68, x75_c, x76, x79, x80_c, x84, x85, x88, x91_c, x93);
and (w5140, x0, x1_c, x2_c, x3_c, x4_c, x6_c, x8, x9_c, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17_c, x20_c, x21_c, x22, x23, x24, x25, x27, x28_c, x29_c, x30_c, x31_c, x32_c, x33, x34, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x43_c, x44, x45_c, x48, x49_c, x50, x51_c, x53_c, x54, x55_c, x56, x58_c, x59, x60, x61, x62_c, x63, x64, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x71, x73_c, x74, x75, x76_c, x78, x79_c, x80, x81, x82_c, x85, x86_c, x87_c, x88, x89_c, x90_c, x91, x93, x94, x95_c, x96_c, x97_c, x98_c, x99);
and (w5141, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5142, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14, x16, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5143, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5144, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5145, x0, x1, x2_c, x3_c, x4, x5, x6, x7_c, x8_c, x9, x10, x11_c, x12, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31, x32, x33_c, x34, x35_c, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43, x44_c, x45_c, x46, x47_c, x48, x49_c, x50_c, x51_c, x52_c, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61, x62_c, x63, x64, x65_c, x66, x67_c, x68_c, x69, x70, x71_c, x72_c, x73, x74, x75_c, x76, x77, x78, x79, x80, x81, x82_c, x83_c, x84, x85_c, x86_c, x87, x88_c, x89_c, x90, x91_c, x92, x93, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w5146, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x72_c, x81, x84, x85, x95, x99);
and (w5147, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30_c, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5148, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5149, x0_c, x2_c, x7_c, x12_c, x24_c, x25, x27, x29_c, x30_c, x31, x35, x38, x40_c, x49, x59, x60, x71_c, x72_c, x73_c, x94, x95);
and (w5150, x0, x1, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5151, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5152, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x85_c, x86_c, x87, x88_c, x89, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5153, x3_c, x4, x8, x10, x14_c, x16, x19_c, x24, x29, x33, x34, x35_c, x38, x42, x43_c, x47_c, x48, x49, x50, x52_c, x53_c, x58, x60, x61_c, x63, x64, x65, x71_c, x74_c, x76_c, x77_c, x80_c, x81, x82, x87, x90, x92_c, x95, x96);
and (w5154, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5155, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5156, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5157, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x25, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5158, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x73_c, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5159, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x37, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5160, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88, x89, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5161, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5162, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62, x82, x90_c, x96, x98, x99_c);
and (w5163, x12_c, x32, x91, x93, x94_c, x95, x96, x97_c, x98, x99);
and (w5164, x0_c, x1, x2, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5165, x8, x21_c, x25_c, x27_c, x34, x39, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5166, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x62_c, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5167, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89, x90_c, x92, x94_c, x95_c, x96_c, x97_c, x99_c);
and (w5168, x5_c, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5169, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91, x92, x93_c, x94, x95_c, x96, x98_c);
and (w5170, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5171, x5, x9_c, x11_c, x12_c, x14, x18, x20, x26, x30, x32, x33, x35, x42, x44, x45, x47, x48_c, x51_c, x53_c, x55_c, x58, x59, x66_c, x70, x71_c, x73_c, x74_c, x75_c, x80_c, x82, x83_c, x86_c, x94, x98_c);
and (w5172, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x67, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5173, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5174, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73_c, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w5175, x2_c, x3_c, x4, x5, x7_c, x8, x9_c, x10, x11_c, x12_c, x14, x15, x16, x17, x18, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27_c, x28, x29_c, x30, x32, x33_c, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x42_c, x43, x44_c, x46, x47_c, x48, x49, x50, x53, x54, x55, x56_c, x57_c, x59_c, x60_c, x63_c, x64_c, x65_c, x66, x67, x68, x69, x70_c, x71_c, x73_c, x75_c, x76, x77_c, x78, x79, x80_c, x81_c, x82_c, x83, x84, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94, x95_c, x96, x97, x98);
and (w5176, x2_c, x3_c, x4, x5_c, x6_c, x7, x8_c, x9_c, x11_c, x12_c, x13, x15_c, x16_c, x17, x18, x19, x20, x22, x23, x24_c, x25, x27, x29, x30, x31_c, x34, x35, x36_c, x37, x39, x40, x41, x42, x43_c, x44, x45_c, x46, x48_c, x49_c, x50, x51_c, x52, x54, x55, x57, x58, x59_c, x61, x62, x65, x66, x67_c, x68, x69, x70, x72, x73_c, x74, x75_c, x77_c, x79_c, x80, x81, x82_c, x83, x84, x86, x88_c, x90, x91, x92, x93_c, x94_c, x95, x98, x99);
and (w5177, x0, x2, x4_c, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5178, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5179, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x53_c, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5180, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5181, x4_c, x6, x7, x8, x9, x11, x13_c, x14_c, x15, x16_c, x18_c, x20, x21_c, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34_c, x35, x36_c, x37, x39, x40, x41, x42_c, x43, x47_c, x48, x49, x50_c, x52, x53_c, x54_c, x55, x56, x58, x59_c, x61_c, x63, x65_c, x67, x68_c, x69_c, x70, x71, x72_c, x74, x75, x76_c, x77_c, x79_c, x80, x82_c, x83_c, x84_c, x86_c, x90, x91, x93_c, x95, x98);
and (w5182, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5183, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w5184, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42, x71_c);
and (w5185, x0_c, x2, x3_c, x5, x7, x9_c, x11, x13, x16_c, x19_c, x22, x23_c, x24_c, x27_c, x28_c, x31_c, x32, x36_c, x38, x43, x49_c, x50_c, x52_c, x53, x56_c, x58, x59_c, x62_c, x64, x65, x66_c, x67_c, x68_c, x72_c, x73, x78, x83, x84_c, x88, x91, x93, x96, x97, x98_c, x99_c);
and (w5186, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x93_c, x94_c, x95_c, x97_c);
and (w5187, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34_c, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5188, x0, x1_c, x2_c, x3, x4_c, x5_c, x6_c, x8, x9, x10, x11, x12, x13, x14_c, x15, x16, x17, x18_c, x19_c, x20, x21, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33_c, x34, x35_c, x36, x37, x38_c, x39_c, x40, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51_c, x52, x53, x54, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62_c, x63_c, x64, x65, x66, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78, x79_c, x80, x81_c, x82_c, x83_c, x85, x86_c, x87_c, x88_c, x89_c, x90_c, x91, x92, x93, x94_c, x95, x96_c, x97, x98_c, x99_c);
and (w5189, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5190, x0, x4_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5191, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5192, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x74_c, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5193, x2, x9, x11, x15, x16, x17_c, x18_c, x19_c, x23, x24_c, x25, x27_c, x28_c, x29, x30, x35, x36_c, x39, x40_c, x41_c, x44_c, x47, x48_c, x51, x55_c, x58, x68, x70_c, x73_c, x74_c, x75, x76, x77_c, x78, x81, x82_c, x83_c, x86_c, x88, x89_c, x95, x96_c, x97_c);
and (w5194, x8, x21_c, x25_c, x27_c, x34, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5195, x11, x12_c, x15, x17_c, x19_c, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5196, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x65_c, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5197, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5198, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5199, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91_c, x92, x93, x94_c, x95, x98, x99_c);
and (w5200, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w5201, x2_c, x4_c, x8, x9, x11_c, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5202, x12_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5203, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5204, x12_c, x40, x74_c, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5205, x0_c, x1_c, x2_c, x4_c, x5_c, x6_c, x7_c, x8, x9, x10, x11, x12, x13, x14, x15, x18, x23, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34, x35, x39, x40_c, x42_c, x44, x45_c, x47, x49_c, x50, x53_c, x54, x55_c, x57, x58, x59_c, x60, x62_c, x63_c, x67_c, x68, x70, x71_c, x73, x74_c, x76, x77, x78, x80_c, x81, x86, x87_c, x88_c, x89_c, x90, x91, x93_c, x95, x96, x97_c, x98);
and (w5206, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x83_c, x93_c, x97_c);
and (w5207, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x65_c, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w5208, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x79, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5209, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x75, x84_c, x85_c, x97_c);
and (w5210, x0_c, x2, x3, x5, x6, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19_c, x20, x21, x22, x23, x25, x28_c, x29, x30, x31, x32, x33, x34_c, x35_c, x36_c, x37, x38, x39, x40, x41_c, x42_c, x43_c, x44, x46_c, x47_c, x48, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57_c, x58, x59, x60, x61, x62, x63_c, x64, x65, x66, x67_c, x68_c, x69_c, x71, x72_c, x73_c, x74_c, x75, x76_c, x78_c, x79_c, x80, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91_c, x93_c, x94_c, x96, x97_c, x98, x99);
and (w5211, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55, x82, x90_c, x96, x98, x99_c);
and (w5212, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5213, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5214, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60_c, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5215, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x90, x93, x97_c, x98_c, x99_c);
and (w5216, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91, x92, x93_c, x94_c, x96, x98, x99);
and (w5217, x49, x83_c, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5218, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5219, x2_c, x11, x23_c, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5220, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92, x93, x94, x96, x97_c);
and (w5221, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5222, x0, x1_c, x2_c, x3, x4, x5, x6, x7, x10, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5223, x4_c, x5_c, x7_c, x8, x9, x83_c);
and (w5224, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5225, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x16, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5226, x13_c, x14_c, x24, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w5227, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x35_c, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5228, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52_c, x71_c);
and (w5229, x0, x1, x2, x5, x7, x9_c, x11, x12, x13_c, x14, x16, x17, x18, x19, x20, x21, x22_c, x24, x26_c, x29, x30_c, x31_c, x32_c, x33, x34, x36, x37, x38, x40_c, x41_c, x43, x46_c, x47_c, x48, x49, x50, x51, x52, x55_c, x57, x59_c, x60_c, x61, x65_c, x66, x69_c, x70_c, x71_c, x72, x73, x74_c, x78_c, x80, x81_c, x83_c, x84_c, x86, x88, x89, x90, x91_c, x93_c, x94, x95_c, x97_c, x99_c);
and (w5230, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x32, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5231, x0_c, x1_c, x2_c, x3_c, x4_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x15, x16_c, x17, x18_c, x19_c, x20_c, x21, x22, x23, x24, x25, x26, x28_c, x30, x31, x32_c, x33, x34, x35, x36, x37, x38, x39_c, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48_c, x49_c, x50, x51, x52, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x63, x64, x65, x66, x67_c, x70, x71, x73_c, x74, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x83, x85, x86, x87, x88_c, x89_c, x90_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99_c);
and (w5232, x0, x1, x3, x4, x5, x6_c, x7, x8, x9, x10, x11_c, x12_c, x13_c, x14_c, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23_c, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40, x41, x42_c, x43, x44, x45_c, x46, x47, x48, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57, x58, x59, x60, x61_c, x62, x63, x64, x65_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85, x86_c, x87, x88, x89_c, x90, x91, x92_c, x93, x94, x95_c, x96, x97_c, x98, x99_c);
and (w5233, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x59, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5234, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x26, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5235, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88_c, x93_c, x97_c);
and (w5236, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x68, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5237, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5238, x11, x12_c, x15, x17_c, x19, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5239, x0, x1, x2, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w5240, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5241, x0, x2_c, x4, x10, x12, x13_c, x16, x23_c, x24, x25_c, x32, x33_c, x35, x36_c, x41, x49_c, x50_c, x53_c, x56_c, x62, x63_c, x65_c, x67_c, x74_c, x75_c, x82, x84_c, x87, x88_c, x92, x93, x94_c, x97);
and (w5242, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x73, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5243, x8, x9_c, x16, x24, x25, x26, x32_c, x40, x42_c, x45, x48, x60_c, x63, x69_c, x87, x91, x94, x98_c, x99_c);
and (w5244, x0_c, x1, x2_c, x4, x7, x9_c, x12_c, x13, x15_c, x16, x17, x18, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x31, x32, x34, x36, x39_c, x40, x41, x42_c, x44_c, x45_c, x46_c, x49_c, x50_c, x51_c, x52, x53, x54, x55, x57_c, x58_c, x61_c, x62, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x73, x76_c, x77_c, x81_c, x82, x83, x86, x88, x89, x90, x91_c, x93, x94, x95_c, x96_c, x97, x98, x99);
and (w5245, x12_c, x40, x65, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5246, x2, x3_c, x4, x6_c, x8, x10, x12_c, x13_c, x16, x19, x21, x22_c, x23_c, x25, x26_c, x28, x29_c, x30, x31_c, x34, x35, x36_c, x39, x41, x42_c, x43_c, x44_c, x45_c, x50, x51, x52, x55, x59_c, x61_c, x62_c, x64, x65_c, x67_c, x68_c, x70_c, x71, x72, x73_c, x74, x75, x76, x77_c, x79, x80_c, x81, x82_c, x83, x86, x87, x88, x89, x91, x92, x93, x94_c, x97, x99);
and (w5247, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5248, x1_c, x4_c, x8_c, x9_c, x10, x13_c, x14_c, x18, x23, x30_c, x33, x38, x39, x40, x42, x44_c, x50, x51_c, x56_c, x57, x58_c, x76, x84_c, x91, x94, x95_c, x98, x99);
and (w5249, x0, x1_c, x3_c, x4_c, x6, x7, x8_c, x10_c, x11, x12_c, x13, x14, x15, x16, x17_c, x18, x19_c, x20, x21, x22, x24, x25_c, x26_c, x27, x28, x30, x31, x32, x34_c, x36_c, x37_c, x38_c, x39_c, x40, x41_c, x42_c, x44, x45, x46, x47_c, x48, x50_c, x51_c, x52_c, x53, x54_c, x56_c, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75, x76_c, x79_c, x80_c, x81_c, x82, x83, x84, x85_c, x86, x87_c, x88_c, x89_c, x91, x92_c, x94_c, x95_c, x96, x97_c, x99);
and (w5250, x71_c, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5251, x16_c, x18_c, x19_c, x20, x22, x26, x32_c, x35, x40, x44_c, x46, x47, x53, x55, x58, x61_c, x64, x65, x68, x71_c, x72, x75, x78, x81_c, x83, x89_c, x90, x94_c, x95_c, x98);
and (w5252, x0, x1_c, x2, x3, x5_c, x6, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5253, x1_c, x3, x7, x8, x9_c, x10, x11_c, x13_c, x14_c, x15_c, x16, x17_c, x18, x20, x21_c, x24_c, x25, x28_c, x30, x36_c, x37, x41, x44_c, x48, x54, x58, x59, x62_c, x66_c, x68, x69, x71_c, x72, x73_c, x80_c, x82, x86_c, x87, x95);
and (w5254, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x30_c, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5255, x0, x1, x2, x4_c, x6_c, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5256, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x60_c, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5257, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x35_c, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5258, x0, x1, x2_c, x3, x4, x5_c, x6, x7, x8, x9_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29, x30, x31_c, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x39_c, x40, x42_c, x43, x44, x45_c, x46, x47, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x56, x57, x58_c, x59_c, x60, x61_c, x62, x63, x64_c, x65_c, x66_c, x67, x68, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x77_c, x78, x79, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x89_c, x90, x91, x93_c, x94_c, x95_c, x96, x97, x98);
and (w5259, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x64_c, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5260, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5261, x1_c, x3, x4, x8, x9_c, x11, x13_c, x14_c, x15_c, x16, x17, x23_c, x24_c, x29_c, x30, x31_c, x35_c, x38_c, x39_c, x40, x44, x45_c, x46, x49_c, x52_c, x53, x56_c, x62, x64, x65_c, x66, x68, x72_c, x73_c, x76_c, x78, x79_c, x81_c, x83_c, x84, x86_c, x87, x88_c, x89, x90_c, x91, x92_c, x99);
and (w5262, x1_c, x2, x5, x6, x8_c, x9, x10_c, x15, x16_c, x23_c, x27, x28, x29, x31_c, x40, x41_c, x43_c, x44, x46, x48_c, x52, x53, x54, x56_c, x57, x60_c, x61, x62, x63, x67, x68, x82_c, x88_c, x90_c, x92, x93_c, x98_c);
and (w5263, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89, x90_c, x92, x94_c, x95_c, x96_c, x98, x99_c);
and (w5264, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w5265, x0_c, x1, x2_c, x3, x4_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5266, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5267, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76, x81, x84, x85, x95, x99);
and (w5268, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x90_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5269, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5270, x1_c, x3_c, x4, x5, x7_c, x8, x9, x11_c, x13_c, x14, x16_c, x17, x18, x20, x21, x22_c, x26_c, x27_c, x28, x35, x38_c, x39, x41_c, x52_c, x57, x59_c, x72_c, x74_c, x77_c, x78, x80, x85_c, x88, x93_c, x98);
and (w5271, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97_c, x98, x99);
and (w5272, x30, x36, x40_c, x55, x60_c, x63, x67, x73, x95_c);
and (w5273, x0, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5274, x0, x1_c, x2_c, x3, x4_c, x5_c, x6, x8_c, x9_c, x10_c, x11, x12, x14, x15, x16, x17_c, x18_c, x19, x20_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x30, x31_c, x32_c, x33_c, x34, x36_c, x37_c, x38_c, x40_c, x41, x42_c, x43, x44_c, x45, x46, x47_c, x48, x49, x50_c, x51_c, x52_c, x53_c, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62, x64, x65_c, x66_c, x67, x68_c, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x75, x77, x78, x79, x80, x81_c, x82_c, x83, x84, x85_c, x86_c, x87, x88, x89, x90_c, x91, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w5275, x15, x24, x33, x37_c, x56_c, x65_c, x82, x94, x98);
and (w5276, x0_c, x1_c, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5277, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5278, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5279, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x43_c, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5280, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5281, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89_c, x97_c);
and (w5282, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x95_c, x97_c, x99_c);
and (w5283, x21, x30, x39_c, x50_c, x54_c, x64, x71_c);
and (w5284, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x64, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5285, x56, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5286, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5287, x5, x9_c, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5288, x0, x1, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5289, x0, x3, x10, x13, x14, x15, x16_c, x22, x24, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5290, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w5291, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5292, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5293, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x95, x96_c, x97_c, x98, x99_c);
and (w5294, x7, x22, x29, x36, x37_c, x40_c, x41_c, x44, x47, x48_c, x49_c, x53, x56_c, x67_c, x68_c, x78_c, x79, x84, x89_c, x90_c);
and (w5295, x5, x10, x16, x20, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w5296, x12_c, x27, x63, x70, x80_c, x88_c, x89, x93);
and (w5297, x0_c, x1, x2, x4_c, x5_c, x6_c, x8_c, x9_c, x10, x11, x12, x13_c, x14, x15, x16_c, x17_c, x18, x19, x20_c, x21, x22, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35_c, x37_c, x38, x39_c, x40, x41_c, x43, x44_c, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52, x53, x55, x56_c, x57, x58_c, x59, x60_c, x61, x62_c, x63, x64_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71_c, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83, x84, x85, x86, x87, x88_c, x89_c, x90_c, x91_c, x92, x93_c, x94_c, x95_c, x96_c, x97, x98, x99_c);
and (w5298, x0_c, x4_c, x5_c, x6_c, x8_c, x10, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5299, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x45_c, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w5300, x26_c, x29_c, x31, x36_c, x38_c, x39, x47, x56, x63_c, x68_c, x78, x84_c, x86, x88_c, x89_c, x92, x93, x97);
and (w5301, x8, x21_c, x25_c, x27_c, x33, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5302, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x89, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5303, x0_c, x1, x2, x3_c, x4_c, x5, x7, x10, x11_c, x13_c, x15, x18_c, x19_c, x21_c, x23_c, x27_c, x28, x29_c, x30_c, x34, x36_c, x37, x38_c, x40_c, x41_c, x42, x45_c, x47, x48, x49_c, x50, x52_c, x54_c, x56_c, x57_c, x58_c, x62, x63, x65_c, x66_c, x67, x68, x71_c, x74, x75, x77_c, x78, x79, x80_c, x81, x82_c, x88_c, x91, x94, x95_c, x96_c, x98_c, x99_c);
and (w5304, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x84_c, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5305, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5306, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5307, x0, x3, x10, x13, x14, x15, x16_c, x17_c, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5308, x0_c, x1_c, x2, x4, x5_c, x6, x7, x8_c, x9_c, x10, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x19, x20, x21, x22, x24, x27_c, x28, x29_c, x30_c, x31, x32, x33, x35_c, x36_c, x37, x38_c, x39, x40_c, x41, x44_c, x46_c, x47, x48_c, x49_c, x51, x53_c, x54_c, x55, x56_c, x60, x61_c, x62, x63_c, x66_c, x67, x68, x69_c, x70, x71_c, x72, x73, x75, x76, x77_c, x78_c, x79, x80, x81, x82, x83_c, x84, x85_c, x86, x87, x88_c, x89_c, x92, x93_c, x94_c, x95, x96, x97_c, x98_c);
and (w5309, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x57_c, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5310, x0, x3_c, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5311, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5312, x0_c, x1_c, x2_c, x3, x4_c, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13, x14_c, x15_c, x16, x17, x18_c, x19_c, x20, x21, x22_c, x23, x24_c, x25_c, x26, x27_c, x28_c, x29, x30_c, x31_c, x33_c, x34_c, x35_c, x36_c, x37_c, x38, x39_c, x41_c, x42, x43_c, x44, x46_c, x47, x48_c, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56, x57_c, x58_c, x59, x60_c, x61_c, x62, x63_c, x64_c, x65, x66_c, x67, x68, x69, x70_c, x72_c, x73, x74, x75, x76, x77, x78_c, x79_c, x80_c, x82_c, x83, x84_c, x85_c, x86_c, x87, x88, x90_c, x91, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5313, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5314, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5315, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89_c);
and (w5316, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5317, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97_c, x98, x99);
and (w5318, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5319, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x59_c, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5320, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80_c, x90_c, x93_c, x97_c);
and (w5321, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x71_c, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5322, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5323, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x50_c, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w5324, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x66_c, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5325, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5326, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5327, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x67, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5328, x0_c, x2, x3_c, x5_c, x6, x7, x10_c, x14_c, x15_c, x17, x20_c, x21, x22_c, x23_c, x24_c, x27, x28_c, x29, x30_c, x31, x34, x36_c, x37_c, x38, x39_c, x41_c, x43_c, x44_c, x46_c, x50_c, x51, x52, x54, x55_c, x57_c, x58_c, x59, x62_c, x63, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x82, x83, x84, x86_c, x87, x88, x89_c, x90_c, x91_c, x92, x94_c, x95_c, x96, x99_c);
and (w5329, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x36_c, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5330, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5331, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5332, x13_c, x14_c, x37_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5333, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5334, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5335, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x73, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5336, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x54, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5337, x0, x4, x5, x6, x8, x9, x11, x12, x13, x15_c, x16, x17, x18_c, x19, x23_c, x24_c, x26_c, x27, x28_c, x29_c, x31, x35, x37, x38_c, x39_c, x40, x41, x42_c, x43_c, x44_c, x49_c, x52, x53_c, x54, x56, x57_c, x62, x63_c, x65_c, x66_c, x69, x70, x72_c, x74, x76, x78, x79, x80, x83_c, x85, x86_c, x88_c, x91_c, x92, x95_c, x96_c, x97_c, x98);
and (w5338, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x82, x90_c, x96, x98, x99_c);
and (w5339, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x44_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5340, x8_c, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5341, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38_c, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5342, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w5343, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5344, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x81, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5345, x12_c, x27_c, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5346, x0_c, x5, x23_c, x30, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5347, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5348, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x86_c, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5349, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5350, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5351, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5352, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w5353, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5354, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x53_c, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5355, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x83);
and (w5356, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5357, x33, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5358, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w5359, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5360, x0, x1, x2_c, x3, x4, x5_c, x6_c, x8_c, x10_c, x12, x13_c, x14, x15, x16_c, x17, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27_c, x28_c, x29_c, x30_c, x31_c, x32_c, x33, x34, x35_c, x37_c, x38, x40, x41, x42_c, x43, x44_c, x46_c, x48, x49_c, x50, x51_c, x52, x53_c, x55, x56, x57, x59, x60_c, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x68_c, x69_c, x70_c, x71_c, x72, x73_c, x74_c, x75, x76_c, x78, x79, x80, x81_c, x82_c, x83_c, x84_c, x86, x87, x88_c, x90_c, x92_c, x95, x96, x97_c, x99_c);
and (w5361, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x97, x98_c, x99_c);
and (w5362, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5363, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x54_c, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5364, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x82, x88_c, x93_c, x95_c);
and (w5365, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5366, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x87, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5367, x11_c, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5368, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x12, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5369, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5370, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5371, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5372, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x48, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5373, x14, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5374, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x96_c, x98, x99_c);
and (w5375, x0_c, x1, x2_c, x5, x10, x11_c, x13, x16_c, x17, x19, x22, x24, x25_c, x26_c, x32, x33_c, x38, x40_c, x41, x42_c, x46_c, x47, x49, x51, x52_c, x53, x56_c, x58_c, x59, x62, x63, x64_c, x66_c, x69, x70, x72, x73_c, x76, x77, x84_c, x86_c, x90_c, x94_c, x95, x96_c, x97_c, x99);
and (w5376, x3, x4_c, x9, x15_c, x16_c, x19_c, x20_c, x21_c, x22_c, x24, x27_c, x33, x37_c, x43_c, x44, x58_c, x63_c, x67, x72_c, x77_c, x80_c, x84, x90_c, x93, x99);
and (w5377, x12_c, x14);
and (w5378, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5379, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x69, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5380, x8, x20_c, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5381, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5382, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x15, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5383, x0_c, x1_c, x5_c, x6, x7, x8, x10_c, x11_c, x12, x13_c, x17, x18, x19, x20, x21_c, x26, x27, x30, x31, x32, x33, x35_c, x36, x37, x38_c, x39_c, x40_c, x41, x43_c, x44, x46, x48, x49, x50, x51, x52, x55, x56_c, x57, x58_c, x60, x62, x63, x64_c, x65, x66, x67, x69, x70_c, x71, x72_c, x73, x76, x78_c, x81, x82, x83_c, x84_c, x85, x86, x87_c, x88_c, x90_c, x91, x92_c, x94_c, x95, x96, x97);
and (w5384, x0, x26_c, x30_c, x36_c, x37, x48, x74_c, x96);
and (w5385, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x89_c, x91_c, x92, x93, x94_c, x97_c);
and (w5386, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x74_c, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5387, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5388, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x86, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5389, x6, x9_c, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5390, x1, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5391, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54_c, x83_c);
and (w5392, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x49, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5393, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x54, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5394, x0_c, x5, x16_c, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5395, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5396, x0_c, x2_c, x4, x5, x7, x8_c, x9, x10_c, x12, x13_c, x20_c, x21, x24, x25, x29, x31_c, x32, x33, x34, x35, x36, x37_c, x38, x45, x49, x50_c, x54, x55_c, x56, x58_c, x59, x62_c, x63_c, x65_c, x73_c, x75_c, x77, x79, x80_c, x81, x83, x86_c, x90_c, x91_c, x92_c, x93, x94_c, x97_c, x98, x99_c);
and (w5397, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x75_c, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5398, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5399, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5400, x0_c, x5_c, x6, x7, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5401, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39, x40, x82, x90_c, x96, x98, x99_c);
and (w5402, x0_c, x1, x2, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x11, x12, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21, x22, x23, x24_c, x25_c, x26, x27, x28_c, x29_c, x30, x31_c, x32_c, x33, x34_c, x35, x36_c, x37_c, x38_c, x39_c, x40, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50_c, x51_c, x52_c, x53_c, x54, x55, x56, x57, x58, x59, x60, x61_c, x62, x63, x64, x65, x66_c, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85_c, x86, x87, x88_c, x89, x90, x91, x92, x93, x94_c, x95_c, x96_c, x97, x98, x99_c);
and (w5403, x8, x16, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5404, x7_c, x9_c, x13, x14, x21, x45_c, x50_c, x59, x61_c, x63_c, x65_c, x72, x77_c, x78, x79, x83, x84, x89_c);
and (w5405, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5406, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5407, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x53, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5408, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20, x40, x82, x90_c, x96, x98, x99_c);
and (w5409, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x93, x95_c, x96_c, x97_c);
and (w5410, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5411, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5412, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5413, x0_c, x1, x2, x3, x4, x5, x6, x7, x8_c, x9, x10_c, x11, x12, x14, x15, x16, x17_c, x18, x19, x21_c, x22, x23, x24_c, x25_c, x26, x27_c, x28_c, x31, x32_c, x33, x34, x35, x36, x37_c, x38, x40_c, x41_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x52, x53_c, x56_c, x57, x58, x59_c, x60, x61_c, x62_c, x63, x64, x66_c, x67_c, x68_c, x70, x71_c, x72, x73, x75, x78, x79_c, x81, x82_c, x83, x84, x85_c, x86, x88_c, x89_c, x90_c, x91_c, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w5414, x8_c, x11_c, x12_c, x14, x15_c, x19_c, x24, x26_c, x28_c, x32_c, x33_c, x39_c, x40, x47, x48_c, x57_c, x66, x69, x70, x76, x77_c, x91_c, x95_c, x98);
and (w5415, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5416, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5417, x0, x1, x2, x5, x6_c, x7, x12, x14, x15, x16_c, x17_c, x19, x22_c, x23, x25, x26, x27, x29_c, x30, x31_c, x32, x33, x34_c, x36_c, x39, x40_c, x41_c, x44, x45_c, x47_c, x48_c, x49, x51_c, x52_c, x54, x56, x57, x58_c, x59_c, x60_c, x61_c, x62_c, x66, x67_c, x68_c, x70, x71_c, x72, x73_c, x74_c, x76_c, x78, x79, x80, x81_c, x82_c, x83, x85_c, x86, x87_c, x88, x90, x91_c, x92, x93_c, x94_c, x97_c, x98, x99);
and (w5418, x0, x2, x3_c, x6_c, x8_c, x9, x10_c, x11, x13_c, x15, x16, x17, x18_c, x19_c, x20_c, x21, x24_c, x25_c, x26, x27_c, x28, x29, x30, x32, x33, x34, x35_c, x38_c, x40, x41, x44, x45, x46, x47, x48_c, x50, x51, x53_c, x55_c, x57_c, x59_c, x60_c, x61_c, x62_c, x63_c, x64, x68_c, x69, x70_c, x71_c, x72_c, x73, x74, x76_c, x77_c, x81, x82_c, x83, x84, x85, x87_c, x89_c, x90_c, x91_c, x93, x97, x99);
and (w5419, x5_c, x9, x27_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5420, x0, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5421, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x13, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5422, x3_c, x4_c, x5_c, x6_c, x7_c, x9_c, x11, x13, x15, x22_c, x23, x24_c, x25_c, x28, x31_c, x32, x34_c, x36_c, x40_c, x42_c, x43_c, x46_c, x49, x53_c, x54_c, x55, x58_c, x59_c, x72_c, x75_c, x76_c, x79_c, x80, x82_c, x84_c, x94, x99_c);
and (w5423, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5424, x0_c, x2_c, x6_c, x7, x8_c, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w5425, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x53, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5426, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x39_c, x40_c, x41_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5427, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53_c, x83_c);
and (w5428, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5429, x11_c, x15_c, x16, x18, x21, x28, x71_c);
and (w5430, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x8, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5431, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5432, x12_c, x23, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5433, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x67, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5434, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x85_c, x89, x93, x97_c, x98_c, x99_c);
and (w5435, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x85_c, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5436, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x30_c, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5437, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78_c, x82, x90_c, x96, x98, x99_c);
and (w5438, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x41, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5439, x0_c, x2, x3, x4, x5_c, x9_c, x12_c, x13, x15_c, x16_c, x17_c, x18_c, x21, x22, x23, x25_c, x27, x28, x29, x30_c, x33_c, x34_c, x35, x39_c, x41, x43, x45_c, x46_c, x47, x50_c, x52, x53, x54_c, x55, x61_c, x63, x64_c, x65_c, x67, x68, x69, x71_c, x72, x76_c, x77_c, x79, x81, x82, x83, x84_c, x88, x89, x91, x92_c, x95_c, x96, x97, x98, x99);
and (w5440, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x81_c, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5441, x0_c, x2, x3_c, x8_c, x12, x22, x24_c, x28_c, x29_c, x33, x35, x39, x40_c, x46_c, x48, x53_c, x55_c, x60_c, x66, x72, x75_c, x78, x82, x83, x86, x87, x95, x96_c, x97_c);
and (w5442, x0_c, x1, x2_c, x3_c, x4, x6, x8, x13, x16, x17, x19, x20, x22, x24, x25_c, x26_c, x27_c, x29_c, x31, x32, x33, x34_c, x35_c, x37_c, x38_c, x39_c, x40_c, x43, x44, x45, x46_c, x47_c, x49, x52, x53_c, x54_c, x55, x56_c, x58, x61, x63_c, x64, x67, x68, x70, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x84_c, x85_c, x88, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x97, x98_c);
and (w5443, x1, x5, x7_c, x17, x18, x19, x20_c, x22, x23, x24_c, x31_c, x32, x35_c, x38, x40_c, x41, x43, x47_c, x49_c, x53_c, x54_c, x57, x58_c, x59, x76, x79_c, x80_c, x81_c, x85, x89_c, x90_c, x91, x99);
and (w5444, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5445, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x38_c, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5446, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5447, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x93_c, x97_c);
and (w5448, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5449, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x83_c, x93_c, x97_c);
and (w5450, x73, x84_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5451, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36_c, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5452, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x98, x99_c);
and (w5453, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w5454, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91_c, x93, x97_c, x98_c, x99_c);
and (w5455, x1_c, x2, x4_c, x11, x12_c, x15, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5456, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74, x75, x84_c, x85_c, x97_c);
and (w5457, x12_c, x32, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5458, x0, x1, x4, x5_c, x6, x7, x8_c, x9_c, x10, x11_c, x12_c, x13, x15_c, x16, x17, x18, x19_c, x20, x21, x22_c, x23_c, x24_c, x25, x27_c, x29_c, x30_c, x31, x32, x33, x35_c, x36_c, x38, x40_c, x41, x42, x43, x45, x46_c, x47, x48, x49, x50_c, x51, x54, x55, x56_c, x57_c, x59_c, x60_c, x61, x62_c, x63, x64_c, x65, x66, x67, x69_c, x70, x72, x73_c, x75_c, x77, x78_c, x79, x81, x82, x83_c, x84, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93_c, x95, x97_c, x98);
and (w5459, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w5460, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5461, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5462, x20_c, x25, x31, x35, x51_c, x68);
and (w5463, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5464, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5465, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x89, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5466, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5467, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46_c, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5468, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5469, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x71, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5470, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5471, x1_c, x9_c, x11_c, x15_c, x28_c, x47, x48_c, x49_c, x56_c, x59, x62, x64_c, x75, x78);
and (w5472, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5473, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5474, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x48_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5475, x12_c, x32, x91, x94, x95, x96, x97_c, x98, x99);
and (w5476, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x69_c, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5477, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94, x97_c);
and (w5478, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5479, x6, x17_c, x20_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5480, x5, x10, x16, x21_c, x30_c, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5481, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29, x40, x82, x90_c, x96, x98, x99_c);
and (w5482, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5483, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5484, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5485, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5486, x0_c, x4, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5487, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x43_c, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5488, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5489, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5490, x0, x1_c, x6_c, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5491, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x77, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5492, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x65, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5493, x3_c, x11, x15_c, x19_c, x20_c, x21, x24_c, x25, x26_c, x31, x33_c, x34, x36, x44, x49, x57, x62, x64_c, x65, x72, x73, x76_c, x78_c, x85, x88, x89_c, x91_c, x93);
and (w5494, x50, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5495, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5496, x2, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5497, x0, x2_c, x6_c, x8_c, x9_c, x10_c, x11_c, x13, x16_c, x19, x20_c, x23_c, x24_c, x25_c, x26_c, x29_c, x30, x31, x33, x36, x39_c, x40_c, x41, x48_c, x50_c, x53_c, x56_c, x57_c, x58, x59, x60, x61_c, x64_c, x65, x71, x77, x78_c, x81, x83, x86, x87, x89_c, x90, x91, x93, x96_c, x98, x99);
and (w5498, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x92, x93, x95_c);
and (w5499, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x58, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5500, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x93_c, x95_c, x96, x98, x99);
and (w5501, x5, x6_c, x13, x14_c, x18_c, x22, x29, x31_c, x34_c, x40_c, x47_c, x53_c, x59, x63, x70_c, x72_c, x73, x77, x78_c, x90_c, x96_c);
and (w5502, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5503, x0, x2, x3_c, x9_c, x14, x15, x21, x25, x26_c, x28, x29_c, x31, x33_c, x35_c, x38, x41_c, x46, x55_c, x63_c, x65, x70_c, x91, x93_c, x95_c);
and (w5504, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5505, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x58, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5506, x8, x17, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5507, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x80, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5508, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5509, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x34, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5510, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x45_c, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5511, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5512, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5513, x5_c, x9, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5514, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x82_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5515, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x87, x88, x91_c, x93_c, x97_c);
and (w5516, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5517, x0_c, x1_c, x2, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5518, x5_c, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5519, x21, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5520, x1_c, x3, x4_c, x6, x7, x8_c, x10, x11_c, x12_c, x13, x15, x16, x18_c, x20_c, x21, x22, x23_c, x25, x26_c, x28, x34_c, x38, x40_c, x42_c, x43_c, x45_c, x46, x49_c, x53_c, x54, x56_c, x60_c, x61, x62, x63, x66, x67_c, x68, x69, x70_c, x72, x73, x75, x76, x78, x79_c, x82, x85, x86_c, x87, x91, x93, x94, x96, x99_c);
and (w5521, x2_c, x3, x4_c, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5522, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5523, x26_c, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5524, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x58_c, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5525, x0, x1, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w5526, x3, x4_c, x6_c, x12_c, x16_c, x23_c, x24_c, x29_c, x31_c, x36_c, x39_c, x45_c, x46, x50_c, x53, x54, x55_c, x56, x62, x68, x70_c, x72_c, x81_c, x83, x89_c, x91, x92_c, x93_c, x96, x97_c);
and (w5527, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5528, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x46, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5529, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5530, x0, x1_c, x2_c, x4, x10_c, x16_c, x17, x18_c, x19, x22, x24_c, x27, x31_c, x32, x35, x36_c, x39, x45, x46, x47_c, x50, x53_c, x54, x59_c, x60, x61, x64, x66_c, x72, x74, x78_c, x86, x91_c, x92_c, x95, x97_c);
and (w5531, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89, x91_c, x92_c, x94, x95_c, x97, x99_c);
and (w5532, x0_c, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5533, x0_c, x5, x23, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5534, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5535, x0, x1_c, x2_c, x3, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5536, x6_c, x8, x12_c, x17_c, x24_c, x26_c, x36, x37_c, x42_c, x43, x48, x49_c, x51, x71, x73_c, x75_c, x76, x80, x95_c, x99);
and (w5537, x0_c, x6_c, x10_c, x11, x13_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5538, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w5539, x2_c, x4, x6, x9_c, x10, x18_c, x29, x30_c, x32_c, x38, x39_c, x40, x44, x52, x53_c, x54, x55, x57_c, x61_c, x62_c, x66, x70_c, x73, x75_c, x76_c, x87_c, x88_c, x91, x99);
and (w5540, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67, x83_c);
and (w5541, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x70, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5542, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x24, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5543, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x59, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5544, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5545, x0_c, x2, x3_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5546, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5547, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x89, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5548, x0_c, x2_c, x4_c, x7, x8, x9, x11, x12, x16, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5549, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5550, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5551, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x92_c, x93, x95, x97_c);
and (w5552, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5553, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5554, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x82_c, x83, x93_c, x97_c);
and (w5555, x0_c, x1, x9, x10_c, x20, x23, x31_c, x35, x39_c, x42_c, x44_c, x47, x50_c, x62, x65_c, x73_c, x76, x77, x79, x81, x83_c, x84_c, x87_c, x91, x99);
and (w5556, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5557, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x97, x99_c);
and (w5558, x5_c, x9, x21, x22, x23_c, x25_c, x26_c, x28_c, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5559, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5560, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5561, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5562, x0_c, x1, x2_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5563, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w5564, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5565, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57_c, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5566, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5567, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5568, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5569, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x52_c, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5570, x38, x39, x84_c);
and (w5571, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62_c, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5572, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5573, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90, x93_c, x97_c);
and (w5574, x1, x5_c, x10, x12_c, x17, x18_c, x19, x26_c, x31, x37, x44, x53, x54_c, x58_c, x62, x63, x65, x68, x72_c, x73, x74, x75, x84_c, x85, x87, x88, x91_c, x94, x95, x96_c);
and (w5575, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w5576, x47_c, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5577, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5578, x2_c, x10, x15, x24_c, x26_c, x27, x28, x35_c, x39, x46, x48, x50, x51_c, x58_c, x61_c, x64_c, x66_c, x69_c, x73_c, x74_c, x76, x81_c, x82, x84, x86_c, x88, x89, x98, x99_c);
and (w5579, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w5580, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x61, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5581, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5582, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x89, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5583, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5584, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5585, x0, x2, x3, x6_c, x10_c, x11, x13_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5586, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x47, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5587, x0, x1_c, x2, x3, x4, x6, x7_c, x8_c, x9, x10_c, x12, x13, x14, x16_c, x17, x18_c, x19_c, x20_c, x21, x22_c, x23, x24_c, x26, x27, x28_c, x29_c, x30, x31_c, x32, x33_c, x36_c, x37, x38_c, x41, x42, x43_c, x44, x46, x47, x48_c, x49_c, x50, x51, x52, x53_c, x54_c, x55_c, x58_c, x59_c, x60_c, x62_c, x64, x65_c, x67_c, x68, x70_c, x71, x72, x73, x74_c, x75, x76_c, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x88, x89, x90, x91, x93_c, x95_c, x96, x97, x99);
and (w5588, x1, x2_c, x5_c, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5589, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52_c, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5590, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5591, x0, x1_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5592, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x82, x83, x93_c, x97_c);
and (w5593, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5594, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5595, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73_c, x79, x90_c, x93_c, x97_c);
and (w5596, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x27_c, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5597, x2_c, x8_c, x25_c, x27, x36_c, x45_c, x47, x62, x72, x73, x75_c, x91, x99_c);
and (w5598, x0_c, x5, x23_c, x27, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5599, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x81, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5600, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5601, x12_c, x40, x82, x87, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5602, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x51_c, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5603, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x56_c, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5604, x2_c, x11, x29_c, x42_c, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5605, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5606, x0, x2, x3_c, x4, x5_c, x7, x8, x9, x13_c, x18_c, x20, x27_c, x29, x30_c, x31, x34, x36_c, x40_c, x42, x43, x47_c, x50, x51, x53, x54, x55, x57_c, x59, x62, x65_c, x66, x71, x75, x77_c, x79_c, x80_c, x81_c, x82_c, x83_c, x84, x87_c, x89);
and (w5607, x0, x1_c, x2, x3, x4_c, x5_c, x6, x7, x11_c, x12, x13, x14_c, x15_c, x16, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36, x38, x39, x40_c, x41, x42, x43, x44_c, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55_c, x56, x57_c, x58_c, x59_c, x60_c, x61, x62_c, x63, x64_c, x65_c, x66, x67_c, x68, x69_c, x70, x71, x72_c, x73_c, x74, x75, x76_c, x77_c, x78_c, x79, x80, x81, x82, x83, x84, x85, x86_c, x87_c, x88, x89_c, x90_c, x91, x92_c, x93_c, x94_c, x95, x96, x97, x99_c);
and (w5608, x0, x2, x3_c, x4_c, x5_c, x8, x9_c, x10, x11_c, x12, x14_c, x15, x16, x17, x18_c, x19, x20_c, x21, x22_c, x23, x24, x25_c, x26_c, x27, x28_c, x29, x30, x33_c, x34, x37, x38_c, x41_c, x43, x44, x45, x46, x47, x48, x51, x52_c, x53, x54_c, x56, x57, x60_c, x61_c, x62, x63_c, x64_c, x65_c, x70_c, x71_c, x73_c, x76, x77, x82_c, x83_c, x84, x85_c, x86, x87, x92_c, x94, x95_c, x96_c, x97, x99_c);
and (w5609, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5610, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69_c, x83_c);
and (w5611, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5612, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x63, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5613, x5, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5614, x14_c, x28, x30_c, x31, x35, x42, x46_c, x53, x54, x55, x76_c);
and (w5615, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5616, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5617, x2, x4, x18_c, x26_c, x30_c, x33, x39, x55_c, x57, x59_c, x66_c, x72_c, x74_c, x88, x92, x94_c, x95, x99);
and (w5618, x49, x72, x73_c, x74, x75, x76, x79, x90_c, x93_c, x97_c);
and (w5619, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5620, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5621, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x83_c);
and (w5622, x0_c, x4_c, x7, x8, x11, x12, x14, x18_c, x21, x25, x30_c, x31_c, x38, x41, x43_c, x44_c, x45, x50, x52, x55_c, x58, x60_c, x68_c, x69_c, x70_c, x71_c, x74, x76_c, x77, x85, x89_c, x90, x93_c, x99_c);
and (w5623, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5624, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5625, x0_c, x1, x2, x3, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5626, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5627, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x82_c, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5628, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64_c, x83_c);
and (w5629, x6_c, x8, x17_c, x26_c, x37, x44, x47_c, x62, x69);
and (w5630, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5631, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x78_c, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5632, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5633, x12_c, x40, x57_c, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5634, x0_c, x1_c, x3, x4_c, x5, x7_c, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5635, x7_c, x26, x35_c, x40, x46_c, x53, x62, x66_c, x68_c, x71, x88_c, x92_c);
and (w5636, x0, x4_c, x6_c, x7_c, x8, x11, x14, x17, x18_c, x19_c, x20_c, x21, x22_c, x24, x25_c, x26, x27, x29, x31_c, x32, x33_c, x35, x36, x38, x39_c, x40, x41_c, x42, x46, x47_c, x48_c, x49_c, x50, x53, x54, x55, x56_c, x57, x58, x59, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68, x70_c, x73, x74, x75, x76_c, x78, x81, x83_c, x85_c, x88_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x98_c, x99_c);
and (w5637, x1, x7, x20_c, x24, x25, x29_c, x44, x56, x71, x91_c, x94, x96_c, x98_c);
and (w5638, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x95, x97, x98, x99_c);
and (w5639, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68, x83_c);
and (w5640, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5641, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5642, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5643, x37, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5644, x3, x13, x24, x27_c, x29, x31_c, x33_c, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5645, x12_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5646, x8, x11_c, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5647, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5648, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5649, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5650, x5, x10_c, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w5651, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5652, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x47, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5653, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x34, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5654, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5655, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5656, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91_c, x92, x93, x94, x95_c, x96, x98, x99);
and (w5657, x2_c, x11, x29_c, x52, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5658, x49, x70, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5659, x1_c, x2_c, x4_c, x7, x19, x22, x23, x28_c, x30_c, x33_c, x38, x43_c, x44_c, x52, x64, x72, x74, x76, x79_c, x82, x89_c, x94_c, x95, x99_c);
and (w5660, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5661, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5662, x0_c, x3_c, x4_c, x6_c, x8_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5663, x0, x1_c, x2_c, x3, x5, x6_c, x7, x8_c, x9_c, x10_c, x11_c, x13_c, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x21, x23_c, x24, x25_c, x26, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34, x35, x36_c, x37_c, x38, x39, x40_c, x41, x42_c, x43, x44_c, x45_c, x46, x47_c, x48, x49, x50_c, x51, x52, x53, x54, x55, x56, x57, x58_c, x59, x60, x61, x62, x63, x64, x65_c, x67, x68, x69_c, x70_c, x72_c, x73_c, x75_c, x77, x78_c, x80_c, x81, x82, x83, x84, x85, x86, x87_c, x88_c, x90_c, x91, x92, x93, x94, x95_c, x97, x98, x99_c);
and (w5664, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x93_c, x97_c);
and (w5665, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76_c, x77, x82, x83, x93_c, x97_c);
and (w5666, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89, x90_c, x94_c, x95_c, x97_c);
and (w5667, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x31, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5668, x0, x4_c, x9_c, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5669, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5670, x13_c, x14_c, x37_c, x39, x40, x82, x90_c, x96, x98, x99_c);
and (w5671, x2, x8_c, x10, x14, x16, x22_c, x23, x24, x27, x29_c, x31, x32, x33, x36, x38_c, x40, x42_c, x45_c, x46_c, x50, x59, x63, x68_c, x76, x85_c, x87_c, x89, x91, x95, x97_c, x98_c);
and (w5672, x45, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5673, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w5674, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23_c, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5675, x0, x2, x4, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x22_c, x24_c, x25_c, x26, x29, x30_c, x33, x34, x35_c, x36_c, x37_c, x40_c, x41_c, x46_c, x48, x51, x52_c, x53_c, x54_c, x55_c, x57_c, x59, x60_c, x64_c, x65, x68_c, x70_c, x71_c, x72_c, x73_c, x74, x77, x78, x79_c, x81, x82_c, x83_c, x84, x85, x87_c, x89, x91, x92_c, x97, x98, x99_c);
and (w5676, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x39, x40_c, x41_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5677, x22, x34_c, x55, x63_c, x76_c, x80, x91);
and (w5678, x0, x3, x4, x5, x8, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5679, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64, x65, x72_c, x81, x84, x85, x95, x99);
and (w5680, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69, x75, x84_c, x85_c, x97_c);
and (w5681, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97, x98, x99_c);
and (w5682, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5683, x0, x1_c, x2_c, x4, x5_c, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5684, x7_c, x8, x15_c, x18_c, x19, x20, x23_c, x25_c, x36, x44_c, x51_c, x57, x59_c, x62, x64_c, x70, x74, x79, x80, x81_c, x90_c, x91_c, x97_c, x99_c);
and (w5685, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94, x95, x99);
and (w5686, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5687, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5688, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5689, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x8_c, x9_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w5690, x6, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5691, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96, x97_c);
and (w5692, x12_c, x40, x82, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5693, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5694, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5695, x18, x42_c, x45, x51, x58);
and (w5696, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5697, x0, x1, x2, x3, x4, x5, x6, x7_c, x8, x9, x10_c, x12, x13, x15, x16, x17, x18, x19_c, x20_c, x21_c, x22, x23_c, x25_c, x26, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x41_c, x42_c, x43, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51_c, x52_c, x53_c, x54, x55, x56_c, x57, x58_c, x59, x60, x61_c, x62_c, x63, x64_c, x65, x66, x67_c, x68_c, x69, x70, x71, x72_c, x73, x74_c, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97, x98_c, x99_c);
and (w5698, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x58, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5699, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5700, x1_c, x3_c, x7, x8, x9, x10, x11_c, x12_c, x13_c, x14, x18, x20_c, x21, x25_c, x26, x27_c, x28_c, x29, x30, x33, x38, x43, x44, x45_c, x48, x50_c, x51, x52_c, x53_c, x55, x58, x61_c, x62_c, x63_c, x64_c, x66_c, x67, x68, x70_c, x71, x72, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x82_c, x84, x85_c, x87, x89_c, x92_c, x93_c, x94_c, x95, x97, x99);
and (w5701, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w5702, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x68, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5703, x1, x8_c, x13_c, x14, x15_c, x16_c, x17, x18_c, x20, x22, x23_c, x24_c, x25_c, x26_c, x27, x29, x30, x32_c, x33, x34, x36, x37_c, x38, x40_c, x54, x58_c, x59_c, x60, x61, x62_c, x63, x64_c, x65_c, x66, x68_c, x69, x70, x71, x73, x76_c, x77, x79, x81_c, x82, x83_c, x84, x85, x90, x92, x93_c, x96, x99_c);
and (w5704, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5705, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x57_c, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5706, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x63, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5707, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5708, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92, x93_c, x95_c, x96, x98, x99);
and (w5709, x49, x63, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5710, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99_c);
and (w5711, x0, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5712, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x95_c, x96_c, x97, x98, x99_c);
and (w5713, x0_c, x1_c, x2_c, x3, x4, x6, x7, x8, x9_c, x10, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17, x18, x19, x20_c, x21, x22_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x38_c, x39_c, x40_c, x42, x44, x45, x46_c, x49, x51_c, x52_c, x53, x54, x55, x57, x58_c, x59, x60_c, x61, x62, x63, x64, x66, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x75_c, x76, x77_c, x78_c, x80, x81_c, x82_c, x83_c, x84_c, x85, x86, x87_c, x88, x89, x90, x91, x93, x94_c, x95, x96_c, x97, x98_c, x99_c);
and (w5714, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x90_c, x92_c, x94, x95_c, x96, x97, x99_c);
and (w5715, x3, x11, x27, x34_c, x40_c);
and (w5716, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5717, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x62, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5718, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x19, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5719, x0, x1_c, x2_c, x3_c, x5_c, x6, x7, x8_c, x9, x10_c, x11, x12, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24, x25, x26, x27, x28, x29_c, x30, x31, x32_c, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x54, x55_c, x56_c, x58_c, x59_c, x60, x61, x63_c, x64, x65, x66, x67, x68, x69_c, x70, x71_c, x72, x73, x74, x75, x76, x77, x78_c, x79, x80, x81_c, x82_c, x83_c, x84, x85_c, x86, x87, x88, x89, x90_c, x91_c, x92, x93_c, x94, x95, x96, x97_c, x98_c, x99_c);
and (w5720, x0_c, x1_c, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11_c, x12_c, x13, x14, x15_c, x16, x17, x18, x19_c, x20, x21, x22, x23_c, x24_c, x25, x26_c, x27_c, x28, x29, x30_c, x31, x32, x33, x34_c, x35_c, x36_c, x37, x38_c, x39, x40, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52_c, x53, x54, x55_c, x56_c, x57_c, x58_c, x59, x60_c, x61, x62_c, x63, x64, x65, x66, x67, x68, x69, x70, x71_c, x72_c, x73_c, x74, x75_c, x77_c, x78_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90, x91_c, x92, x93_c, x94, x95_c, x96, x97_c, x98_c, x99);
and (w5721, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x16, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5722, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5723, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5724, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5725, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x26_c, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5726, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77, x84_c, x85_c, x97_c);
and (w5727, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5728, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39_c, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w5729, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x65, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5730, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5731, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5732, x8, x21_c, x25_c, x27_c, x34, x39_c, x42, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5733, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5734, x0, x6_c, x7_c, x14, x16, x19_c, x22_c, x25_c, x29, x33_c, x34_c, x36, x37_c, x39, x42_c, x44, x47, x49_c, x57, x58_c, x59, x61, x62, x67_c, x70, x71_c, x72, x75_c, x78, x79_c, x83, x86, x90_c, x91_c, x95, x98_c);
and (w5735, x0_c, x1, x2_c, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5736, x4, x7, x8, x13_c, x15_c, x19_c, x20, x25_c, x27_c, x30, x35_c, x42, x43_c, x45, x46, x52, x56, x60, x61_c, x62_c, x70, x74_c, x75_c, x83, x87_c, x92_c, x94_c);
and (w5737, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5738, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x56_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5739, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x62_c, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5740, x2_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5741, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x96, x98, x99_c);
and (w5742, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x93, x97_c);
and (w5743, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83_c, x90_c, x96, x98, x99_c);
and (w5744, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x43_c, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5745, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5746, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x21_c, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5747, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5748, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x88, x90_c, x91, x92, x95, x97_c);
and (w5749, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5750, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5751, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x85, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5752, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19_c, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w5753, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5754, x15_c, x19, x23_c, x35_c, x60, x84, x88_c);
and (w5755, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5756, x0, x2, x3, x6_c, x10_c, x11, x13_c, x18_c, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5757, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5758, x0_c, x5, x23_c, x25, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5759, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5760, x0_c, x2_c, x3_c, x7_c, x16, x38_c, x40_c, x42_c, x51, x72, x90, x93, x97);
and (w5761, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80, x85, x89, x93, x97_c);
and (w5762, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x44, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w5763, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5764, x1_c, x2, x4_c, x6_c, x7, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14, x17, x21, x22_c, x24_c, x26_c, x28, x29_c, x32_c, x33, x34_c, x35, x37_c, x38, x39, x42, x43_c, x44, x45, x49, x50, x51_c, x53_c, x54_c, x55_c, x58, x59_c, x60_c, x61_c, x62, x63_c, x64, x65, x66, x67_c, x68_c, x70, x71, x72_c, x73, x74_c, x75_c, x76, x78, x80, x81_c, x82, x83_c, x85, x86, x88_c, x89_c, x95, x96_c, x98_c, x99);
and (w5765, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w5766, x0, x1, x2, x3, x4_c, x5, x8_c, x9_c, x10_c, x11_c, x12, x13, x14_c, x15, x16_c, x17_c, x18, x19_c, x20_c, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32, x33, x34, x35, x36_c, x38_c, x39, x40_c, x41, x42, x44, x45_c, x46, x47, x48, x49, x52_c, x53_c, x55, x57_c, x59_c, x61_c, x62, x63, x64_c, x65_c, x66_c, x69_c, x70, x71, x72_c, x74, x75, x76_c, x77, x79, x81, x82, x83_c, x84, x86_c, x87, x88_c, x89_c, x91_c, x92, x94_c, x95_c, x96, x97_c, x98, x99_c);
and (w5767, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5768, x1, x2_c, x3_c, x6_c, x7, x8, x9_c, x10, x11_c, x12, x15_c, x16, x17, x18_c, x22, x25_c, x26, x34, x35_c, x36_c, x37, x39, x40, x41_c, x42, x47, x48, x49, x51_c, x61_c, x68_c, x69, x71, x72, x74_c, x75, x78_c, x79_c, x88_c, x91_c, x92_c, x93, x94, x95, x96, x97, x98_c, x99);
and (w5769, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5770, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5771, x0, x1, x2_c, x3, x8_c, x9, x13, x14, x15_c, x16, x17_c, x18_c, x20, x22, x23, x25_c, x28_c, x29_c, x30_c, x31, x34, x35_c, x37_c, x38, x40_c, x42, x44, x45_c, x47, x49_c, x50_c, x53, x56, x58, x59, x60_c, x61_c, x62, x66_c, x67, x68_c, x71_c, x73_c, x74, x75_c, x76_c, x77, x79, x81_c, x82_c, x83_c, x84_c, x85_c, x87, x91_c, x92, x94, x95, x96_c, x98_c, x99);
and (w5772, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5773, x0_c, x1, x2, x3_c, x4_c, x5_c, x7_c, x8, x10_c, x11_c, x12_c, x13, x14_c, x16_c, x17_c, x18_c, x20_c, x21, x22_c, x24, x26, x27_c, x28_c, x29_c, x30, x31_c, x32_c, x34, x35_c, x36_c, x39_c, x40, x41, x42_c, x43, x44, x46, x47, x48_c, x49_c, x50, x51_c, x53_c, x54_c, x56_c, x57, x58, x59, x60_c, x62, x63_c, x65, x66_c, x67, x68_c, x69, x70, x71, x73_c, x74, x75, x76, x77_c, x78, x79, x80, x81_c, x82, x85_c, x88, x90_c, x91, x93, x95, x96, x97_c, x98_c);
and (w5774, x0_c, x1, x2_c, x3_c, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5775, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5776, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x32, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5777, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x53_c, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5778, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5779, x0_c, x4_c, x5_c, x6_c, x8_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5780, x0, x1_c, x2, x3, x4_c, x6_c, x7, x8_c, x9, x10, x11_c, x12, x13, x14_c, x15_c, x16_c, x17, x18, x19, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34, x35, x37, x38, x40, x41, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x53, x54_c, x55_c, x56_c, x59_c, x61, x63, x64, x65, x67_c, x68, x69, x72_c, x73, x74, x75_c, x76_c, x78, x79, x80, x81, x82, x83, x85, x86_c, x87, x88, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96_c, x97, x98_c, x99);
and (w5781, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w5782, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x80_c, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5783, x12_c, x40, x62, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5784, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x50, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5785, x13_c, x14_c, x16_c, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w5786, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5787, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5788, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x97_c);
and (w5789, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x76_c, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5790, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x72, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5791, x5_c, x9, x27, x52, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5792, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x66, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5793, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x90_c, x93_c, x97_c);
and (w5794, x19_c, x23, x29_c, x37, x40, x44_c, x45_c, x51_c, x65, x67, x73, x95_c, x97_c);
and (w5795, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x77_c, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5796, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5797, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5798, x0_c, x2, x3, x4, x5_c, x6, x7_c, x8, x9_c, x10, x11_c, x13, x14, x15_c, x16, x17_c, x18, x19_c, x20_c, x21, x22, x23, x24_c, x25, x26_c, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x36, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x44, x45_c, x46, x47_c, x48_c, x49_c, x50, x51, x52, x53, x54_c, x55, x56, x59, x60, x63, x64, x65, x66, x67_c, x68_c, x69, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5799, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89, x90_c, x94, x97_c);
and (w5800, x12_c, x40, x67_c, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5801, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x78_c, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5802, x13, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5803, x0_c, x1_c, x3_c, x4_c, x5, x6_c, x8_c, x9_c, x10_c, x11_c, x13, x14, x15, x16, x17_c, x19, x20_c, x21, x22_c, x23, x24_c, x25_c, x26_c, x28_c, x29, x30, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x39, x40_c, x41_c, x42_c, x43, x44, x46, x47, x48, x50, x51_c, x52, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x61, x62_c, x63_c, x64, x65_c, x66_c, x67_c, x71_c, x72, x73_c, x75_c, x77, x78_c, x79, x80_c, x81, x82, x83, x84, x86, x87_c, x89, x90_c, x92, x93_c, x94_c, x95, x97_c, x98, x99_c);
and (w5804, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5805, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5806, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x82, x83, x93_c, x97_c);
and (w5807, x0_c, x1, x2_c, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5808, x10_c, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5809, x12_c, x24, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5810, x0_c, x2_c, x4_c, x7_c, x9_c, x10_c, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5811, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5812, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5813, x4_c, x6_c, x8, x10_c, x11, x13, x16_c, x18, x19_c, x22, x23_c, x24_c, x35, x38_c, x39_c, x41_c, x43, x46, x48, x49_c, x50, x54_c, x58_c, x63_c, x64_c, x68_c, x70, x73, x74_c, x76, x78_c, x80_c, x81_c, x84_c, x85, x87, x93_c, x95_c, x97_c, x98_c);
and (w5814, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5815, x5_c, x10_c, x20_c, x32, x35, x36, x38, x40_c, x45, x46_c, x47_c, x51, x52_c, x63_c, x66, x73, x77, x79, x90, x91, x93);
and (w5816, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5817, x8_c, x11, x19, x43_c, x44_c, x50_c, x69, x81_c);
and (w5818, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5819, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22, x83_c);
and (w5820, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5821, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x87_c, x93_c, x97_c);
and (w5822, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5823, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5824, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5825, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x51_c, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w5826, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5827, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54, x73_c, x76, x85, x89, x93, x97_c);
assign w5828 = x19;
and (w5829, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40, x83_c);
and (w5830, x13_c, x27_c, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w5831, x0_c, x1, x3_c, x4, x5_c, x8, x9_c, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5832, x0_c, x1_c, x5, x8, x10, x11_c, x20_c, x23, x30, x33_c, x35, x36_c, x37_c, x47_c, x48, x60_c, x62_c, x64_c, x69_c, x70, x72_c, x73, x77, x78_c, x79_c, x83_c, x85_c, x86, x90_c, x92);
and (w5833, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5834, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36_c, x71_c);
and (w5835, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x50, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5836, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5837, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5838, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5839, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x37, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5840, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5841, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x96, x97_c, x98, x99_c);
and (w5842, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x30, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5843, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5844, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5845, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5846, x0_c, x4, x12_c, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5847, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x37_c, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5848, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x95_c, x96_c, x98_c);
and (w5849, x4_c, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5850, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5851, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5852, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5853, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x65_c, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5854, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x43_c, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5855, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5856, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5857, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5858, x12_c, x40, x46_c, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5859, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x79, x90_c, x93_c, x97_c);
and (w5860, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x96, x97_c, x98, x99_c);
and (w5861, x12_c, x18, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5862, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x36_c, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5863, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x66, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5864, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5865, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w5866, x60_c, x69_c);
and (w5867, x3_c, x4, x6, x8, x10, x11_c, x12_c, x14_c, x17, x20_c, x21_c, x22_c, x23, x25, x26_c, x27, x30, x31_c, x32, x33, x35_c, x36, x38_c, x40_c, x41, x42, x48, x49, x50, x51_c, x53_c, x58, x59_c, x60, x62, x64, x66_c, x68, x69_c, x71, x73, x74, x76, x78_c, x79, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x87, x88_c, x89, x90_c, x91, x92, x93, x96, x99_c);
and (w5868, x0, x2, x4_c, x5_c, x7_c, x8_c, x10_c, x11, x12, x13, x14, x16, x18, x19_c, x20_c, x22_c, x24, x31_c, x32_c, x33, x34_c, x38, x39_c, x40_c, x42_c, x43, x47_c, x48_c, x49, x51, x52_c, x53_c, x54, x57, x59_c, x60, x63, x64_c, x66_c, x67_c, x68_c, x69, x70_c, x71, x72, x74_c, x76_c, x77, x78, x80, x82, x84_c, x86_c, x87, x88_c, x95, x96_c);
and (w5869, x1_c, x2_c, x4, x7_c, x8, x9, x11, x15, x16_c, x19, x22_c, x26, x28, x30, x31_c, x32_c, x35_c, x39_c, x44, x45, x46, x57, x58, x61_c, x62_c, x65_c, x66, x67, x68_c, x70, x71_c, x73_c, x75_c, x76_c, x78, x81, x82_c, x83_c, x84, x85_c, x87, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95_c, x99_c);
and (w5870, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5871, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5872, x0_c, x1, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17, x18, x19_c, x20, x21, x22, x23, x24, x25, x26_c, x27_c, x29_c, x30, x31_c, x32_c, x33, x34, x35, x36_c, x37_c, x38_c, x39, x40_c, x41_c, x42, x43, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x52, x53, x54_c, x55, x56, x57, x58_c, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x75_c, x76, x77, x78, x79, x80, x81, x82, x83_c, x84_c, x85_c, x86, x87, x88_c, x89_c, x90, x91, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w5873, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5874, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5875, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5876, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5877, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w5878, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x72, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5879, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91, x92, x93_c, x94, x96, x98);
and (w5880, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67, x75, x84_c, x85_c, x97_c);
and (w5881, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x67_c, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5882, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5883, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30_c, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5884, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x16_c, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5885, x5, x10, x16, x21_c, x34_c, x35, x41_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5886, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x96, x98, x99);
and (w5887, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x97_c);
and (w5888, x2_c, x3_c, x11, x17, x20_c, x25_c, x27_c, x30, x39_c, x42, x43, x50_c, x53_c, x74, x79, x87_c, x91, x93);
and (w5889, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5890, x0, x1, x2, x3_c, x4_c, x5_c, x6, x7_c, x8, x9, x10, x11, x12_c, x13, x14, x15, x16, x17, x18, x19_c, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x27, x28, x29, x30_c, x31, x32_c, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45, x46_c, x47, x48_c, x49_c, x50_c, x51, x52, x53_c, x54_c, x55_c, x56, x57, x58, x59_c, x60_c, x61, x62, x63_c, x64_c, x65, x66, x67, x68_c, x69, x70, x71_c, x72, x73_c, x74, x75, x76, x77, x78, x79_c, x80_c, x81, x82, x83, x84, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w5891, x22_c, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w5892, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x64, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5893, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34, x40, x82, x90_c, x96, x98, x99_c);
and (w5894, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5895, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5896, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5897, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5898, x1_c, x3_c, x5, x7, x9, x11_c, x12_c, x13_c, x15_c, x16, x17, x18_c, x19_c, x20_c, x21, x24_c, x26, x27, x30, x31, x33, x36_c, x37_c, x38_c, x39_c, x40_c, x42, x43_c, x45, x48_c, x51, x52, x56_c, x57_c, x58_c, x60, x61_c, x62, x63_c, x64_c, x66, x67_c, x68, x72, x73, x74, x75_c, x76, x77_c, x78_c, x80_c, x81_c, x83, x85, x86, x87, x90_c, x92, x94, x97, x98_c);
and (w5899, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x40, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5900, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92, x95, x98_c, x99_c);
and (w5901, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x69_c, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5902, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x84, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5903, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5904, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20_c, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w5905, x0, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5906, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x58_c, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5907, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62, x63_c, x65, x72_c, x81, x84, x85, x95, x99);
and (w5908, x3_c, x5, x6, x7_c, x8_c, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5909, x10_c, x27_c, x31, x35_c, x37, x62_c, x63_c, x65, x67, x68, x69, x73, x74_c, x85, x89, x95_c, x98_c);
and (w5910, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5911, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x95, x97_c);
and (w5912, x0_c, x1, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5913, x0_c, x4, x7, x8_c, x10_c, x11, x12, x13_c, x14, x15_c, x16, x18, x19, x21_c, x22_c, x25, x26, x27, x29, x30, x31_c, x32, x33_c, x34_c, x35, x37, x46, x48_c, x50_c, x51_c, x52, x53_c, x55_c, x56, x60, x62, x63, x64_c, x65, x66, x67_c, x68, x71, x72, x73, x74_c, x75, x76, x80, x85_c, x88_c, x92_c, x98_c);
and (w5914, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46, x83_c);
and (w5915, x0, x1, x2, x3, x4, x6, x7, x8, x9, x10, x11_c, x12_c, x13, x14_c, x15_c, x16, x18, x19_c, x20_c, x22, x23_c, x24, x25, x26_c, x27, x28, x29, x30, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38_c, x39_c, x40_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49, x50_c, x51_c, x52, x53, x54, x56, x57_c, x58, x60_c, x61_c, x62, x63_c, x64_c, x65_c, x66, x67_c, x68, x69, x70_c, x72, x73_c, x74, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x82, x83_c, x84_c, x85_c, x86_c, x87, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w5916, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5917, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5918, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w5919, x70_c, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5920, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5921, x0, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5922, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5923, x7_c, x22_c, x28_c, x40, x41_c, x43_c, x45, x54_c, x63);
and (w5924, x0_c, x1_c, x2_c, x3_c, x4, x5, x6, x7_c, x8_c, x9_c, x10_c, x12_c, x13, x14_c, x15, x16_c, x17, x18_c, x19_c, x20, x22_c, x23, x24_c, x25, x26, x27_c, x28_c, x29_c, x30, x31, x32_c, x33_c, x34_c, x36, x38_c, x39, x40_c, x41, x42_c, x43, x44, x45_c, x46, x47, x48_c, x50, x51, x52, x53_c, x54_c, x55, x56, x57, x58, x59, x60, x61_c, x62, x64_c, x65_c, x66_c, x67, x69_c, x70_c, x71_c, x72_c, x73, x74_c, x75_c, x76_c, x77_c, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87_c, x88, x89, x90, x91, x92_c, x93_c, x94_c, x95_c, x96_c, x97, x98, x99);
and (w5925, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5926, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5927, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5928, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x90, x93_c, x95_c, x96, x98, x99);
and (w5929, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5930, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5931, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5932, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5933, x12_c, x39, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5934, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58, x82, x90_c, x96, x98, x99_c);
and (w5935, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5936, x0_c, x3_c, x4_c, x6, x7_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5937, x2_c, x3_c, x4_c, x5, x7, x8_c, x9_c, x10, x11_c, x13_c, x14_c, x15_c, x16_c, x17, x18, x19_c, x21_c, x22, x24, x26_c, x28_c, x29, x30, x31_c, x32_c, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x42, x43, x44_c, x45, x46_c, x47, x49_c, x50_c, x51_c, x52, x53_c, x55_c, x56_c, x57_c, x58, x59_c, x60_c, x64, x65, x66, x67_c, x68, x70, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78, x79, x80_c, x81_c, x82, x84, x86_c, x87, x88_c, x90_c, x91, x94_c, x96, x97, x98);
and (w5938, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5939, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5940, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91, x92, x93_c, x94, x95_c, x96, x98, x99);
and (w5941, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5942, x2_c, x3, x6_c, x8, x11_c, x12, x16, x19_c, x27_c, x31, x33_c, x37, x43, x47_c, x50, x51, x60, x63_c, x64, x65_c, x67_c, x68_c, x69, x70_c, x71_c, x72, x75_c, x76, x78, x80, x81_c, x87_c, x90_c, x92, x95_c);
and (w5943, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x16, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5944, x2, x4, x10, x14_c, x19, x22, x24_c, x47, x55_c, x77, x79, x81, x83);
and (w5945, x1, x4, x5, x8_c, x14_c, x16_c, x17, x19, x20_c, x23_c, x24_c, x25_c, x27_c, x30_c, x31_c, x35, x36_c, x37_c, x40, x43, x47_c, x48, x51, x54_c, x57, x58, x59_c, x60, x62_c, x66_c, x67, x70_c, x72_c, x79_c, x84, x92_c, x94, x95, x96, x97, x98_c, x99_c);
and (w5946, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x57_c, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w5947, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98_c);
and (w5948, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89, x90_c, x93, x97_c);
and (w5949, x12_c, x32, x60_c, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5950, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5951, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5952, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5953, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10_c, x11_c, x12, x13, x14, x15_c, x16_c, x17_c, x18, x20_c, x21_c, x22_c, x23_c, x24, x25, x26, x27, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36, x38, x40, x42_c, x43, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x52_c, x53, x54, x55, x56, x57, x58_c, x59, x61_c, x62, x63, x64_c, x65, x66, x67, x69_c, x70, x71, x72, x75_c, x76_c, x77, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90_c, x91_c, x92, x93_c, x94, x95, x98_c, x99_c);
and (w5954, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68_c, x83_c);
and (w5955, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x79, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5956, x8, x21_c, x25_c, x27_c, x28, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5957, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x44, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5958, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5959, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5960, x12_c, x19_c, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5961, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x90_c, x92_c, x94_c, x95, x96, x97, x99_c);
and (w5962, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x30_c, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5963, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x37, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5964, x12_c, x32, x43, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5965, x12_c, x32, x66, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w5966, x1_c, x3, x8, x11_c, x12, x13_c, x15_c, x16, x18, x20_c, x21_c, x23_c, x25_c, x26, x28, x29_c, x31, x33_c, x37_c, x39_c, x40_c, x43_c, x44, x45_c, x46_c, x48_c, x51, x53, x54, x58_c, x59, x62_c, x63, x64_c, x65, x66_c, x69_c, x72, x75_c, x79_c, x80, x83_c, x84_c, x86_c, x96_c, x97, x98_c);
and (w5967, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x66, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w5968, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83, x88_c, x92, x94_c, x95_c, x96, x97_c);
and (w5969, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x57_c, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5970, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w5971, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5972, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x75, x77, x82, x83, x93_c, x97_c);
and (w5973, x0_c, x1_c, x2_c, x10_c, x12, x13_c, x20, x21_c, x22_c, x23_c, x26_c, x28_c, x29, x30, x37, x38_c, x39_c, x41, x44_c, x45_c, x50, x51_c, x52_c, x55, x56_c, x59, x61_c, x62, x63_c, x64_c, x65_c, x68_c, x71_c, x72, x74, x78, x80_c, x82, x83_c, x84, x86_c, x87_c, x91, x99);
and (w5974, x3_c, x8, x12, x19_c, x23_c, x33, x36_c, x42_c, x46_c, x55_c, x56, x59, x61, x64_c, x67, x71, x74, x77, x78_c, x84_c, x88, x93_c);
and (w5975, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w5976, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x41_c, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5977, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5978, x5_c, x9, x27, x61_c, x76, x84, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w5979, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w5980, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x20, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w5981, x3, x5, x6, x7_c, x19, x20, x30_c, x31, x33_c, x34, x36, x40, x43_c, x44, x47_c, x48, x54, x58, x61, x63_c, x66, x67_c, x70_c, x72_c, x76_c, x78, x81_c, x82_c, x83, x84, x89_c, x90, x93_c, x96);
and (w5982, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x81, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5983, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x57, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w5984, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x75, x77, x82, x83, x93_c, x97_c);
and (w5985, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x61_c, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w5986, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75_c, x79, x90_c, x93_c, x97_c);
and (w5987, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x70_c, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5988, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x79, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5989, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x52_c, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w5990, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x84_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5991, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5992, x0, x1_c, x2, x3, x5_c, x6_c, x7, x8_c, x9_c, x10_c, x11, x12, x14, x16_c, x17, x18, x19, x20_c, x21_c, x22_c, x23_c, x25_c, x26_c, x27, x28, x29_c, x30, x31, x32_c, x33, x34, x35_c, x36, x37, x38, x39_c, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x52_c, x53_c, x54, x55_c, x58_c, x59_c, x60, x61, x62, x63, x65, x66_c, x67_c, x69, x70, x71, x72_c, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84, x85, x86, x87, x88, x89_c, x90_c, x91_c, x92, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w5993, x0, x2_c, x3, x4_c, x5, x6, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w5994, x0_c, x3, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x11, x12, x15, x16_c, x17, x18_c, x19_c, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35_c, x36, x37_c, x38, x39, x40, x41_c, x42_c, x43_c, x44, x45_c, x46_c, x48, x49, x50, x51, x52, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64, x65, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x73_c, x74, x75, x76, x77, x78_c, x79, x80_c, x81, x82, x83_c, x84, x87, x89_c, x90_c, x91_c, x92, x93, x94, x95, x96, x97_c, x98, x99_c);
and (w5995, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w5996, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x87, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w5997, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x79, x90_c, x93_c, x95_c, x96, x97, x99_c);
and (w5998, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w5999, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7_c, x8_c, x9, x10_c, x11, x12_c, x13, x15, x16, x17, x18_c, x19, x20_c, x21, x22, x23_c, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30_c, x31_c, x32, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x41, x42_c, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50_c, x51, x52, x53_c, x54, x55, x56_c, x57_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81_c, x82, x83_c, x84, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6000, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6001, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6002, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6003, x8, x17_c, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6004, x12_c, x32, x59, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6005, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x40, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6006, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6007, x1_c, x2, x3_c, x4, x7_c, x9, x11_c, x12_c, x14_c, x15, x19, x20, x22, x24_c, x25_c, x28_c, x31, x32_c, x36, x37_c, x38, x42, x46, x48, x49_c, x52, x54_c, x56_c, x64, x68, x73_c, x76, x77, x79, x81_c, x83, x85, x86, x88, x90_c, x91);
and (w6008, x11, x12_c, x15, x17_c, x23_c, x27, x28_c, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6009, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6010, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85, x90_c, x93_c, x97_c);
and (w6011, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x56_c, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6012, x1, x3, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x12, x13, x14_c, x15, x16, x17_c, x18, x19, x20_c, x22_c, x23_c, x24_c, x25, x26, x27_c, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35, x36, x38, x39, x41, x42, x43_c, x44, x45_c, x46_c, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55_c, x56, x58_c, x60, x61_c, x62, x63, x64_c, x65, x66_c, x68, x69, x70_c, x71_c, x72, x73_c, x74_c, x75, x76, x78, x79_c, x80, x81_c, x82_c, x84, x85_c, x86_c, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94_c, x96, x98_c, x99_c);
and (w6013, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x93_c, x97_c);
and (w6014, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6015, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6016, x1, x3_c, x4_c, x5_c, x6_c, x7_c, x8, x9, x10_c, x11, x12, x13, x14, x15, x16_c, x18, x19, x21, x22, x23, x24_c, x26_c, x27_c, x29, x30_c, x31_c, x32_c, x33, x34, x35_c, x36_c, x37, x38_c, x40, x41, x42, x43_c, x44_c, x45, x46_c, x48, x49_c, x50_c, x52, x53, x54, x55, x56_c, x57_c, x58_c, x59, x60, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x70_c, x71, x72, x73, x75_c, x76, x77_c, x78, x79, x80_c, x81, x82_c, x83, x84_c, x86, x87, x88, x90, x91, x93_c, x94, x95, x96, x97, x98_c);
and (w6017, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6018, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x77_c, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6019, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8, x9, x10_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6020, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x72, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6021, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43, x83_c);
and (w6022, x3_c, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6023, x0, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6024, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w6025, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x98_c, x99_c);
and (w6026, x0_c, x5, x11_c, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6027, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x55, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6028, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x60_c, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w6029, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x98_c, x99);
and (w6030, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x76, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w6031, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88, x90_c, x93_c, x96, x97, x98, x99);
and (w6032, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x99);
and (w6033, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6034, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84);
and (w6035, x0_c, x4_c, x5_c, x6_c, x8_c, x9_c, x12_c, x13, x14_c, x16_c, x17, x18_c, x20_c, x22, x25_c, x26, x27, x29, x30_c, x31_c, x32_c, x36_c, x38, x39_c, x41_c, x43, x44, x45, x48_c, x49, x50_c, x51, x52, x53, x54, x55_c, x56_c, x57_c, x58_c, x60_c, x61, x62, x64, x65, x66, x68, x70, x71, x72_c, x74, x75_c, x76, x77, x78, x79_c, x81_c, x84_c, x85, x88_c, x89, x90, x91_c, x92_c, x97_c, x98_c, x99);
and (w6036, x8, x21_c, x25_c, x27_c, x30, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6037, x73, x82_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6038, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x99_c);
and (w6039, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68_c, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6040, x1, x2_c, x3_c, x4, x6_c, x9, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x22_c, x24_c, x25_c, x27, x28_c, x29, x30_c, x32_c, x35, x38, x39_c, x43_c, x44, x45_c, x47_c, x48, x49_c, x50, x51_c, x52, x53_c, x56_c, x57, x58, x59, x60, x63_c, x65_c, x66_c, x67, x70, x72, x74, x75_c, x78_c, x79, x80, x81_c, x83, x84_c, x85, x88_c, x89, x90_c, x91, x94, x95_c, x97_c, x99_c);
and (w6041, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6042, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x18, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6043, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x47_c, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6044, x2_c, x5_c, x6_c, x7, x8, x9, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6045, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x61_c, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6046, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6047, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6048, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x78_c, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6049, x13_c, x14, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w6050, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x31_c, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6051, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x19_c, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6052, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x57_c, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6053, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x68_c, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6054, x3, x4, x5_c, x6_c, x13_c, x14, x15, x17, x18_c, x20_c, x21, x23_c, x24_c, x25_c, x26_c, x29_c, x32, x35_c, x36_c, x37_c, x39, x41, x45, x46_c, x48_c, x49, x51, x52_c, x53_c, x55_c, x56_c, x57, x59, x62, x63, x64, x65_c, x67, x71, x72_c, x74_c, x76_c, x77_c, x78_c, x79_c, x81_c, x83, x84_c, x85_c, x89_c, x90_c, x92_c, x94, x95, x96_c, x98, x99);
and (w6055, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6056, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x27_c, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6057, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6058, x0_c, x1, x2_c, x3_c, x5, x6, x9, x11_c, x12_c, x13_c, x14_c, x15_c, x18_c, x19_c, x20, x21_c, x24_c, x25, x26, x29, x30_c, x32, x34_c, x35, x36_c, x37_c, x40, x41, x43_c, x44, x48_c, x50_c, x51, x52_c, x53, x56, x57, x60, x62, x64, x66_c, x67_c, x69, x71_c, x72, x74, x75, x76, x80, x86_c, x88, x89_c, x92_c, x98_c, x99_c);
and (w6059, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x37_c, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6060, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27_c, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6061, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31, x40, x82, x90_c, x96, x98, x99_c);
and (w6062, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6063, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47, x49, x64, x71, x72_c, x74_c, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6064, x13_c, x39, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w6065, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6066, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6067, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6068, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x91_c, x93_c, x94_c, x95_c, x96, x98, x99_c);
and (w6069, x0, x4_c, x15_c, x20_c, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6070, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w6071, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76_c, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6072, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32_c, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6073, x2, x10_c, x12_c, x17, x19, x29_c, x31_c, x34_c, x49_c, x50_c, x55_c, x59_c, x72_c, x73, x74, x75, x80, x82, x89_c, x97, x98_c);
and (w6074, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6075, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6076, x5, x10, x12_c, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6077, x2, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6078, x0_c, x2_c, x4, x6_c, x9_c, x10_c, x11, x14_c, x15_c, x16, x21, x23, x25_c, x26_c, x27, x28_c, x29_c, x31, x32_c, x33_c, x36_c, x37, x38, x41_c, x42, x43_c, x44, x45, x46, x49, x50_c, x53_c, x54, x55, x57, x59, x60_c, x65, x69_c, x72_c, x73_c, x79_c, x80, x81_c, x83, x84, x87, x89, x92_c, x93, x94, x95, x96_c, x97_c);
and (w6079, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x93_c, x94_c, x95, x96_c, x98, x99_c);
and (w6080, x0, x2_c, x3, x4_c, x5_c, x7_c, x9_c, x12_c, x13, x14, x15, x17_c, x18, x19_c, x20, x21, x22, x23, x25, x28_c, x29_c, x31, x32_c, x35, x39_c, x40_c, x41, x42, x43, x45, x47_c, x49, x51, x52_c, x54, x55_c, x56_c, x59_c, x60, x62, x63, x64, x65, x66_c, x67_c, x68_c, x69, x71_c, x73_c, x74_c, x75, x76_c, x78_c, x79, x80, x81_c, x84_c, x86, x87_c, x89, x90_c, x92_c, x93, x96_c, x98_c, x99_c);
and (w6081, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x64_c, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6082, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x40, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6083, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15_c, x16, x17_c, x19_c, x20, x21_c, x22, x23_c, x24, x25, x26, x27_c, x29_c, x31_c, x32, x33_c, x35_c, x36, x37, x38, x40, x41_c, x42_c, x43_c, x44, x46_c, x47_c, x48, x50_c, x51, x52, x53, x54, x55, x56, x57, x58_c, x59, x61_c, x62, x63_c, x64, x65, x66_c, x67_c, x68_c, x69_c, x71, x72, x77, x78, x79_c, x80, x81, x82, x83, x84, x87_c, x88, x89_c, x91, x92, x95, x96, x97, x98, x99_c);
and (w6084, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6085, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x22, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6086, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6087, x9_c, x10, x11, x12, x14, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6088, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w6089, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w6090, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w6091, x1_c, x3, x10_c, x11, x12, x15_c, x16_c, x18_c, x20_c, x22, x23_c, x24, x26, x28_c, x29, x35, x36, x39_c, x41, x43_c, x45_c, x46, x48, x49_c, x51, x52_c, x53_c, x56_c, x57_c, x60_c, x61, x64, x67, x68_c, x69_c, x73, x74, x75, x79, x81_c, x85, x86, x90_c, x92_c, x96, x97, x99_c);
and (w6092, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w6093, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x87_c, x89, x93, x94_c, x96, x97);
and (w6094, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x29_c, x31_c, x32, x83_c);
and (w6095, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39_c, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6096, x11, x23_c, x71_c);
and (w6097, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x13_c, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6098, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x81_c, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6099, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w6100, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w6101, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6102, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x90_c, x91, x95, x96, x97, x99_c);
and (w6103, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6104, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x40_c, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6105, x51_c, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6106, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x71);
and (w6107, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w6108, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6109, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x55, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6110, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6111, x9_c, x11_c, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6112, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58_c, x60, x61, x62_c, x75, x82_c, x90_c, x96, x98, x99_c);
and (w6113, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6114, x0_c, x1_c, x2, x3, x4_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22_c, x23_c, x24, x25, x26_c, x27_c, x28_c, x29, x30_c, x31, x32, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58_c, x59_c, x60, x61, x62_c, x63, x64, x65, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80_c, x81, x82, x83, x84_c, x85, x86_c, x87, x88, x89, x90, x91, x92_c, x93, x94_c, x95_c, x96_c, x97, x98_c);
and (w6115, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x30, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w6116, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6117, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6118, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x66, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6119, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6120, x0_c, x2_c, x4, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6121, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x68, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6122, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64, x71_c);
and (w6123, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6124, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6125, x4_c, x10, x15_c, x17, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w6126, x0, x1, x2, x4, x9, x10_c, x11_c, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6127, x10, x15, x16_c, x32, x43_c, x52_c, x54, x55_c, x59_c, x63, x71, x81_c, x85_c);
and (w6128, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97, x98_c, x99_c);
and (w6129, x0_c, x3_c, x4_c, x6, x7_c, x10, x11_c, x12_c, x40, x82, x90_c, x96, x98, x99_c);
and (w6130, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6131, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6132, x9, x10, x16_c, x17_c, x21_c, x25_c, x38_c, x55, x61_c, x63, x83, x89, x96);
and (w6133, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c, x97, x98_c, x99_c);
and (w6134, x9_c, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6135, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x70_c, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6136, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6137, x0_c, x1, x2, x3, x4, x6_c, x7, x8_c, x9_c, x10_c, x11_c, x12, x13_c, x14_c, x15_c, x17, x18, x20_c, x21_c, x22_c, x23, x24, x25_c, x26, x27, x28_c, x29, x30_c, x31, x32, x33, x34, x36, x37, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46_c, x48, x49, x50, x51_c, x52_c, x53, x55_c, x56_c, x57, x58, x59, x61_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x73, x75, x78_c, x80, x81_c, x82, x83_c, x84_c, x85_c, x86_c, x87, x88, x89, x90, x91, x92, x93_c, x94, x96_c, x98, x99);
and (w6138, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x83, x93_c, x97_c);
and (w6139, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6140, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6141, x0, x6_c, x7, x10_c, x11, x12, x13, x15, x18, x19_c, x22_c, x25_c, x26_c, x27, x28_c, x30, x31_c, x33, x34_c, x38, x42_c, x43, x44_c, x46_c, x47_c, x53, x54_c, x55, x56, x57_c, x58, x62_c, x64, x66, x67, x68, x69, x70, x72, x73_c, x74, x75, x81, x83, x85, x89_c, x90, x91_c, x92_c, x96, x98, x99_c);
and (w6142, x0_c, x6, x8_c, x10_c, x11, x12_c, x13_c, x14, x15_c, x16_c, x17, x18_c, x22_c, x23, x28_c, x31, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x41, x43_c, x49, x51, x52_c, x53, x54, x55_c, x57_c, x60, x61_c, x62, x63_c, x66, x67, x70_c, x72, x74, x75, x77_c, x79_c, x80, x82_c, x84, x85, x86, x87_c, x89_c, x96_c, x97);
and (w6143, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x51_c, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6144, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6145, x64_c, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6146, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6147, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60_c, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6148, x6, x17, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6149, x49, x65, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6150, x0, x1, x2_c, x3, x5, x7_c, x8, x9, x10_c, x12_c, x14_c, x15_c, x16_c, x17, x18, x20_c, x21_c, x22, x23_c, x25, x26, x27_c, x28_c, x29, x30, x32, x34_c, x35_c, x36, x37_c, x38_c, x39, x40, x42, x43, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50_c, x51, x52_c, x53_c, x54_c, x56, x57_c, x58_c, x59, x60_c, x62_c, x63, x64, x65, x67, x68, x69_c, x70, x71, x72_c, x73_c, x75, x76, x77_c, x78_c, x79_c, x81_c, x82, x83, x84, x86, x87, x88_c, x89, x90_c, x91_c, x92_c, x93, x95, x96, x97_c, x98);
and (w6151, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x76, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6152, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w6153, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x31_c, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6154, x0, x2, x3, x6_c, x7, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6155, x12_c, x32, x36, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6156, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6157, x2, x5_c, x7, x28_c, x32_c, x33_c, x36, x41_c, x57, x62_c, x73_c, x75, x80_c);
and (w6158, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38_c, x83_c);
and (w6159, x12_c, x32, x65_c, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6160, x0, x2, x4, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6161, x5, x10, x16, x21_c, x34_c, x35, x41_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6162, x1, x4_c, x10_c, x11_c, x13_c, x14, x15_c, x19_c, x22, x24, x25_c, x28_c, x31, x35_c, x36_c, x39_c, x41_c, x45, x50, x54, x62, x63, x64, x66_c, x72_c, x76_c, x77, x82, x87, x90, x96_c, x99_c);
and (w6163, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c, x99);
and (w6164, x0, x1_c, x3, x4_c, x6, x7_c, x8_c, x9_c, x10, x11_c, x12, x13, x14, x15_c, x16, x17_c, x18, x20_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x30, x33, x34_c, x35_c, x38, x43_c, x44, x45, x47, x48, x49, x50_c, x51, x52_c, x53, x54, x55, x58_c, x59, x61, x62_c, x64, x65_c, x67, x69_c, x70_c, x71_c, x73, x74_c, x75_c, x76, x79, x80, x81, x82, x85_c, x86_c, x87_c, x88, x90, x91_c, x92_c, x93_c, x94_c, x95, x97, x98, x99);
and (w6165, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11, x83_c);
and (w6166, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x33, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6167, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x54, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6168, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97, x98, x99);
and (w6169, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6170, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6171, x0, x1, x2, x3_c, x4_c, x5_c, x6, x7, x8_c, x9, x10, x11, x12, x13, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27, x28, x29, x30, x31_c, x32, x33, x34, x35, x36, x37_c, x38_c, x39, x40, x41_c, x42, x43, x44, x45_c, x46, x47, x48, x49_c, x50, x51, x52_c, x53, x54_c, x55_c, x56, x57, x58_c, x59, x60_c, x61, x62, x63_c, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73_c, x74, x75, x76, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91, x92_c, x93, x94_c, x95, x96_c, x97_c, x98, x99);
and (w6172, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6173, x0, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6174, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6175, x0, x3, x10, x13, x14, x15, x16_c, x22, x30_c, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6176, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6177, x4_c, x9, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w6178, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55_c, x82, x90_c, x96, x98, x99_c);
and (w6179, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6180, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88, x89_c, x90, x91_c, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6181, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6182, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x47_c, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6183, x0_c, x1, x2, x3, x4, x5_c, x6, x7, x8, x9, x10_c, x11, x12, x13_c, x15, x16, x17, x18, x19, x20, x21_c, x22, x25_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x33_c, x34_c, x35_c, x36, x37, x39_c, x40, x41_c, x42_c, x43_c, x44, x45_c, x46, x47, x48_c, x49, x51, x53_c, x54, x55_c, x57_c, x58, x59_c, x60_c, x61, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69_c, x70_c, x71, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x80, x81_c, x82, x84_c, x85_c, x86, x87, x88_c, x89_c, x90, x91, x92, x93_c, x95, x97, x98, x99_c);
and (w6184, x3_c, x4_c, x6, x9_c, x10_c, x12_c, x13_c, x19, x20_c, x21_c, x24, x28, x31_c, x32_c, x33_c, x39, x40, x41_c, x42, x45, x47, x56, x57, x60, x62, x63, x69_c, x70, x72, x75_c, x76, x79_c, x81_c, x83, x84, x91_c, x95_c, x96_c, x97);
and (w6185, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31, x83_c);
and (w6186, x8, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6187, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x90_c, x92, x95, x96, x97, x99_c);
and (w6188, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x93, x97_c);
and (w6189, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6190, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x97_c);
and (w6191, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x72, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6192, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6193, x2, x4_c, x5, x6, x7_c, x9_c, x13, x15, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6194, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41_c, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6195, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87_c, x88, x89, x90_c, x91, x92, x95, x97_c);
and (w6196, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x16_c, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6197, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6198, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75_c, x76, x85, x89, x93, x97_c);
and (w6199, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x98_c, x99_c);
and (w6200, x0, x1, x2_c, x3, x5, x6, x7, x8, x9, x10_c, x11, x13, x14_c, x15_c, x16, x17, x18, x20_c, x23, x24_c, x26_c, x28_c, x29_c, x30_c, x31, x32, x33, x35, x36, x37_c, x38_c, x39_c, x40_c, x41, x42_c, x44, x47_c, x48_c, x50, x51, x52, x53_c, x54_c, x55_c, x56, x57_c, x59_c, x61, x62, x64, x65, x66, x68_c, x69, x70_c, x73, x74, x76, x77, x78, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85, x86, x89, x91_c, x92_c, x93_c, x95, x96_c, x97_c, x99_c);
and (w6201, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53, x83_c);
and (w6202, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24, x40, x82, x90_c, x96, x98, x99_c);
and (w6203, x1_c, x2, x4, x5_c, x6, x8, x9_c, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6204, x39_c, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6205, x0, x2_c, x4_c, x8, x9, x11, x12, x16, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6206, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6207, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6208, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6209, x1_c, x4, x5_c, x9, x13, x15_c, x18_c, x19, x21, x22_c, x26_c, x27, x30_c, x31_c, x32_c, x35, x38_c, x40, x46, x48_c, x49, x50, x51_c, x52, x55, x56, x57_c, x60_c, x72, x73, x76, x79, x82_c, x84, x85_c, x87, x88_c, x90_c, x91_c, x94_c, x98_c);
and (w6210, x49, x74_c, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6211, x0, x3_c, x4, x5_c, x6_c, x8_c, x13, x20_c, x28_c, x37_c, x38, x41, x43_c, x44, x45_c, x47_c, x50, x56_c, x58_c, x60, x61, x62, x63, x66_c, x67_c, x72_c, x73, x75, x78_c, x81_c, x85, x87, x88, x97_c);
and (w6212, x0, x1, x2_c, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x11_c, x12, x13, x14_c, x15, x16, x17, x18_c, x19, x20_c, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33_c, x34_c, x35, x36, x37, x38, x39_c, x40, x41, x42, x43, x44_c, x45_c, x46, x47_c, x48, x49_c, x50_c, x51, x52_c, x53, x54_c, x55_c, x56, x57, x58, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66_c, x67_c, x68_c, x69, x70, x71, x72_c, x73, x74, x75_c, x76_c, x77, x78, x79, x80, x81, x82_c, x83_c, x84, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91, x92, x93, x94, x95, x96_c, x97_c, x98_c, x99);
and (w6213, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6214, x5, x10_c, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6215, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6216, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6217, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6218, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6219, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6220, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x74_c, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6221, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x96_c, x97_c, x98, x99_c);
and (w6222, x0, x1, x5_c, x11_c, x14, x26, x31_c, x32_c, x34_c, x35, x36_c, x37_c, x38, x45_c, x51, x52_c, x53_c, x54_c, x62_c, x63, x72_c, x76, x77, x81, x82, x83_c, x85, x86_c, x88_c, x92, x94, x98_c);
and (w6223, x2_c, x3_c, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6224, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6225, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x25, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6226, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6227, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6228, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6229, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x44, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6230, x0_c, x1_c, x2, x3_c, x4, x5, x7, x8_c, x10, x11, x12_c, x13_c, x16_c, x17_c, x19_c, x20_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x28_c, x29, x30, x31, x32, x33_c, x34_c, x35, x36_c, x37_c, x38, x40, x41_c, x43, x44_c, x45_c, x47_c, x48_c, x50_c, x51_c, x53, x54_c, x55_c, x57_c, x58, x59, x61_c, x62_c, x63, x64, x65, x66, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75, x76_c, x77, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84, x85, x86_c, x87, x89, x90, x92, x93, x94, x95, x96_c, x97, x98, x99);
and (w6231, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6232, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x83, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6233, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x15, x16, x17_c, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6234, x5, x10, x16, x21_c, x32_c, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6235, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w6236, x5, x10, x16, x21_c, x34, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w6237, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x67_c, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6238, x0, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6239, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x72_c, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6240, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6241, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6242, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x55, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6243, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6244, x0, x2_c, x4_c, x5_c, x7_c, x9, x11, x13_c, x14_c, x15_c, x17_c, x19, x22, x23, x28_c, x32, x33, x36_c, x37_c, x39, x48_c, x50_c, x53_c, x54, x55, x58_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x67_c, x68, x70_c, x71_c, x78, x79_c, x81, x82_c, x83, x85, x86, x87, x89, x90_c, x91_c, x94_c, x95_c, x97, x98_c, x99);
and (w6245, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w6246, x13_c, x14_c, x18_c, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w6247, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x69, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6248, x6_c, x21_c, x39_c, x55_c, x57_c, x62, x65_c, x67, x72, x75, x95, x96);
and (w6249, x1, x3_c, x4_c, x6, x7, x8, x10_c, x12, x13, x14_c, x16, x18_c, x20_c, x22, x23, x24_c, x26_c, x27, x29, x33, x34_c, x35, x36_c, x39, x41, x42, x43, x46_c, x48, x53, x54, x56, x57, x58, x61, x62_c, x63, x64, x68_c, x71_c, x73, x76_c, x77_c, x78_c, x80, x86_c, x89, x93_c, x99);
and (w6250, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6251, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6252, x0_c, x5, x23_c, x26_c, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6253, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49_c, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6254, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6255, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6256, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6257, x0_c, x2_c, x6, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w6258, x1, x2, x3_c, x4, x5_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13, x14_c, x15, x16_c, x17_c, x18_c, x19, x20, x22_c, x23, x24, x25, x26_c, x27, x28, x29_c, x30_c, x31_c, x33_c, x34, x36, x37, x38_c, x39, x40_c, x41_c, x42, x43_c, x44, x45_c, x46, x47_c, x48, x49_c, x51, x52, x53_c, x54_c, x56, x57_c, x58_c, x59, x60_c, x61_c, x62_c, x63, x64_c, x65, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x73_c, x75_c, x76, x77, x78_c, x79_c, x80, x81, x82_c, x83_c, x84, x85_c, x86_c, x87, x88, x89_c, x90_c, x91, x92_c, x93, x94, x96, x97, x98_c);
and (w6259, x7_c, x11, x19, x20, x21_c, x23, x28_c, x31_c, x35_c, x37, x39, x41_c, x42, x45_c, x47_c, x52, x53, x56_c, x68, x84_c, x90, x91, x92);
and (w6260, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x54_c, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6261, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6262, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30_c, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6263, x12_c, x32, x62, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6264, x1_c, x2_c, x5_c, x6, x7_c, x9_c, x11, x12_c, x16_c, x17_c, x22, x23, x24, x26, x27, x28_c, x31, x32_c, x36, x37, x38_c, x39, x40, x42_c, x44_c, x45_c, x47, x48_c, x49_c, x50, x51, x52_c, x53_c, x54, x56, x57, x59_c, x61, x62, x65, x66, x67_c, x68_c, x70, x71, x74, x77_c, x78_c, x79, x80, x81_c, x83_c, x84, x85, x86_c, x87_c, x89, x90, x91_c, x92_c, x96_c, x99);
and (w6265, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6266, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6267, x14_c, x22, x41_c, x42, x76, x79_c, x87, x95, x96, x98_c);
and (w6268, x8_c, x21_c, x44_c);
and (w6269, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6270, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x18, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w6271, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68, x70, x73, x82, x90_c, x96, x98, x99_c);
and (w6272, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6273, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6274, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x62, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6275, x0, x2, x5_c, x6, x7_c, x8_c, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6276, x73, x96_c, x98, x99);
and (w6277, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49_c, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6278, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6279, x1_c, x5, x10_c, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6280, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6281, x11, x12_c, x15, x17_c, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6282, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x99);
and (w6283, x0_c, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6284, x0, x1, x2, x3_c, x5_c, x6_c, x7_c, x8_c, x9, x10, x11_c, x12_c, x14, x15_c, x16_c, x17_c, x18, x19, x20, x21, x22, x23, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31_c, x32_c, x33, x34_c, x35, x36_c, x37_c, x38, x39, x40, x41, x42, x43, x44_c, x45, x46_c, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54, x55_c, x56_c, x57_c, x58_c, x59_c, x60, x61, x62_c, x63, x64_c, x65, x66, x67, x68_c, x69_c, x70, x72_c, x73_c, x74, x75_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99_c);
and (w6285, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x50, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6286, x11, x21, x27, x33_c, x53_c, x60, x72_c, x84_c, x85_c, x87);
and (w6287, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w6288, x0_c, x1, x2_c, x3, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6289, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x39_c, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6290, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6291, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6292, x3_c, x8_c, x18, x27_c, x45, x49_c, x50, x51, x53_c, x56, x68_c, x83_c, x84, x89, x92_c);
and (w6293, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x67, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6294, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x30_c, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6295, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6296, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39_c, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6297, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6298, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6299, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6300, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6301, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6302, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6303, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6304, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6305, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98);
and (w6306, x8_c, x37, x54);
and (w6307, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6308, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6309, x0, x1_c, x2_c, x3, x4_c, x5_c, x6_c, x7_c, x9_c, x10_c, x11, x12_c, x13, x14_c, x15_c, x17_c, x18_c, x19, x20_c, x21, x22, x23, x24_c, x25, x26, x27_c, x28_c, x29, x30_c, x31, x32_c, x33, x34, x35_c, x37_c, x38_c, x39, x40_c, x41_c, x42, x43_c, x44_c, x46, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54, x55_c, x56_c, x57, x58_c, x59, x60_c, x61_c, x62_c, x63, x64, x65, x66, x67_c, x68, x70, x71, x72, x73_c, x74, x75_c, x76, x77_c, x78, x79_c, x80, x81, x82, x83_c, x84, x85, x86_c, x87, x88_c, x89, x90_c, x91_c, x92_c, x93, x95_c, x96_c, x97_c, x98, x99);
and (w6310, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x61, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6311, x10, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6312, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6313, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w6314, x8, x19_c, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6315, x10_c, x21, x34_c, x44, x45_c, x52, x68_c, x69, x73, x78, x82_c, x83, x88, x94, x99);
and (w6316, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6317, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x96, x97_c);
and (w6318, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c, x99_c);
and (w6319, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x40, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6320, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x76, x77_c, x80, x81_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6321, x0, x2_c, x4_c, x6, x7, x9_c, x10, x11, x13_c, x15, x17, x18, x19, x20, x22, x23, x25, x26_c, x28, x29_c, x31_c, x33_c, x35_c, x36_c, x37_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x46, x49_c, x51, x52, x55_c, x58_c, x60, x65_c, x66, x67_c, x69, x70_c, x71, x73, x74, x75, x78, x80_c, x81, x82, x84_c, x86_c, x87, x89, x91, x94, x96_c);
and (w6322, x45, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6323, x0, x2, x7_c, x8_c, x11, x13_c, x15, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6324, x0_c, x4_c, x5_c, x6_c, x8, x12_c, x32, x55, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6325, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6326, x0_c, x5, x8_c, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6327, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6328, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6329, x4_c, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6330, x5, x10, x16, x21_c, x34_c, x35_c, x38_c, x42_c, x46, x47, x50_c, x51, x52_c, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6331, x8, x9_c, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6332, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6333, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x79, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6334, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x30, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6335, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x31_c, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6336, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6337, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6338, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6339, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x77_c, x82, x83, x93_c, x97_c);
and (w6340, x3, x13, x21_c, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6341, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92_c, x94, x95_c, x96, x98, x99);
and (w6342, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15_c, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6343, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x79, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6344, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6345, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6346, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x81_c, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w6347, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x61_c, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6348, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72, x73_c, x76, x85, x89, x93, x97_c);
and (w6349, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6350, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w6351, x6, x15_c, x16_c, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6352, x0, x1_c, x2, x3_c, x4_c, x5, x6, x7, x8, x9, x11_c, x12_c, x13, x14, x15, x16_c, x17, x18, x19_c, x20_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x28_c, x29_c, x30, x32, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x40, x41, x42, x44_c, x45_c, x47, x48_c, x49, x50, x51, x52, x53_c, x54, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x63, x64, x66, x67, x68, x69_c, x70_c, x71_c, x72, x73, x74, x75_c, x76_c, x77, x78_c, x79_c, x80, x81_c, x82_c, x83, x84_c, x85, x86, x87, x88_c, x89_c, x90, x91, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w6353, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x95_c);
and (w6354, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6355, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6356, x0, x41_c, x58_c, x60_c, x63, x83_c, x85);
and (w6357, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6358, x44, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6359, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6360, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6361, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x31_c, x35_c, x39_c, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w6362, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x41_c, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x93, x97_c);
and (w6363, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88, x89_c, x90, x91_c, x92_c, x93, x96_c, x97_c, x98, x99_c);
and (w6364, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6365, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12_c, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6366, x8, x9, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x85, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6367, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x97, x98, x99_c);
and (w6368, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43, x82, x90_c, x96, x98, x99_c);
and (w6369, x8, x21_c, x25_c, x27_c, x34, x37_c, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6370, x0_c, x1_c, x3, x4_c, x5_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6371, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6372, x33_c, x52, x99_c);
and (w6373, x0_c, x5, x21, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6374, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x62_c, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6375, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49, x82, x90_c, x96, x98, x99_c);
and (w6376, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x65, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6377, x5_c, x9, x27, x45, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6378, x20_c, x28_c, x32, x40, x41, x43, x44, x49_c, x52, x55_c, x60_c, x65_c, x71, x72, x73_c, x75, x84, x85_c, x89_c, x92, x93, x98, x99_c);
and (w6379, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x66, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6380, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x66_c, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6381, x0_c, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6382, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6383, x8, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6384, x4_c, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6385, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6386, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6387, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x83_c, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6388, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36_c, x39, x40_c, x41, x44, x46, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6389, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6390, x0_c, x5, x23_c, x24, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6391, x0_c, x3_c, x4_c, x6, x7_c, x10_c, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x93, x95_c);
and (w6392, x0_c, x1_c, x3, x4_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6393, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x39_c, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6394, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x84_c, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w6395, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x66_c, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w6396, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w6397, x21, x22, x23_c, x27_c, x68, x81_c, x83, x94_c, x98);
and (w6398, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93, x95, x97_c);
and (w6399, x0, x2, x6, x7, x8, x9_c, x10, x13_c, x15_c, x16_c, x18_c, x19, x20_c, x22, x25_c, x27, x29, x30, x31_c, x32_c, x34_c, x35_c, x37, x41_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x49, x54_c, x55, x56, x57_c, x62_c, x63, x66, x68, x74_c, x80, x81_c, x82_c, x84, x88_c, x89, x91, x94_c, x99_c);
and (w6400, x0, x3, x4, x5, x8_c, x10, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6401, x0, x2, x3_c, x4, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11, x13_c, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22_c, x23, x24, x25_c, x26_c, x27, x28_c, x30, x31_c, x32_c, x33, x34_c, x35, x36, x37, x38, x39, x40, x41_c, x42_c, x43, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50, x51, x52_c, x53_c, x54_c, x55, x58_c, x59, x61, x62_c, x63_c, x64, x65, x66, x67, x68, x69_c, x70, x71, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78, x79, x80_c, x81, x82_c, x83, x86, x87_c, x88_c, x89, x90, x91_c, x92, x93_c, x94, x95, x96_c, x97_c, x98, x99);
and (w6402, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w6403, x0, x1, x2_c, x3, x4_c, x5, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6404, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6405, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x92, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6406, x6_c, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6407, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6408, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w6409, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6410, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6411, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x40, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6412, x1, x3, x4_c, x5, x7_c, x10_c, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6413, x2_c, x11, x28_c, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6414, x6_c, x9, x29, x66_c, x69_c, x81_c, x82_c, x94_c);
and (w6415, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x76, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6416, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x86, x87, x89, x93_c, x95_c, x96_c, x97_c);
and (w6417, x0_c, x5, x23_c, x30_c, x31_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6418, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6419, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6420, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6421, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x90, x91, x92, x95, x97_c);
and (w6422, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x98, x99);
and (w6423, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92_c, x93, x95_c, x96, x98, x99);
and (w6424, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6425, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6426, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53_c, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6427, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6428, x5, x10, x16, x21_c, x34_c, x35_c, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w6429, x0, x1_c, x2_c, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6430, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6431, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x71, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6432, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x36, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6433, x2_c, x6_c, x9, x10, x11_c, x14, x15, x16, x18, x19, x22, x24_c, x25, x26_c, x27, x28_c, x29, x30, x33_c, x34_c, x35, x36_c, x39_c, x41_c, x42_c, x43, x44, x46, x47_c, x49_c, x50, x52, x54, x55_c, x57, x60, x62, x63, x64, x65_c, x66, x67, x68, x70, x71, x72, x74_c, x75_c, x76, x77, x79, x80, x81, x83, x86, x88, x89_c, x92, x93_c, x94, x95_c, x96_c, x98);
and (w6434, x0_c, x3_c, x4_c, x5_c, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6435, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6436, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19_c, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6437, x0, x2_c, x3, x4_c, x5, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w6438, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x44, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6439, x0, x1_c, x2, x3, x5, x8, x10_c, x11, x12_c, x13, x14, x15, x16, x17, x18_c, x20, x22, x24, x25_c, x27_c, x28_c, x29, x32, x33, x35_c, x38, x40_c, x41, x42_c, x43, x44_c, x47_c, x49, x51_c, x53_c, x54, x56, x58, x59_c, x60, x61_c, x62_c, x63, x64, x69_c, x70, x71, x73_c, x74, x75_c, x77, x78_c, x80, x81, x82_c, x83, x84, x85_c, x86, x87_c, x88, x89_c, x90_c, x94, x97_c, x98, x99);
and (w6440, x12_c, x27, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6441, x0, x2, x7_c, x8, x11_c, x13, x14_c, x27, x28, x30, x53, x55_c, x63, x65, x81, x95, x98_c);
and (w6442, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x18, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6443, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57_c, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6444, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36_c, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6445, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x39, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6446, x8, x11_c, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6447, x3_c, x7, x8_c, x19_c, x30_c, x34, x38_c, x55_c, x61_c, x68, x69, x72, x77, x78, x85_c, x87, x89_c, x94, x95_c, x98);
and (w6448, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17_c, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6449, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6450, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x35_c, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6451, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91, x92, x93_c, x94, x96_c, x98, x99_c);
and (w6452, x2, x4_c, x9_c, x11, x15, x16_c, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6453, x0_c, x3_c, x4_c, x6, x7_c, x8_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6454, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17, x18, x19, x20, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6455, x73, x79, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6456, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53_c, x82, x90_c, x96, x98, x99_c);
and (w6457, x8, x21_c, x25_c, x27_c, x28, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6458, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x24_c, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6459, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6460, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x99);
and (w6461, x4, x9_c, x11, x15, x16_c, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w6462, x4, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27, x40, x82, x90_c, x96, x98, x99_c);
and (w6463, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6464, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6465, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x67, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6466, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6467, x8, x15_c, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6468, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x79, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6469, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x74_c, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6470, x49, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6471, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6472, x23, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6473, x1_c, x5, x9, x11_c, x12, x21, x24, x36, x37, x39_c, x41_c, x42_c, x43_c, x47, x48_c, x53_c, x55, x57, x58_c, x62_c, x67_c, x68_c, x70, x72_c, x74, x76, x77, x84, x85_c, x89, x93_c, x97_c, x98);
and (w6474, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x27, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6475, x12_c, x40, x71_c, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6476, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x49, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6477, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x94_c, x95, x97_c, x99_c);
and (w6478, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x91_c, x93, x95_c, x98, x99);
and (w6479, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31_c, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6480, x12_c, x29, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6481, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x92, x93, x94, x95, x97_c, x99_c);
and (w6482, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86_c, x90_c, x93_c, x97_c);
and (w6483, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6484, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6485, x0_c, x3_c, x5_c, x6, x10, x13_c, x14, x16_c, x17_c, x23_c, x25, x27, x28_c, x29, x31_c, x36, x38_c, x40, x44, x50_c, x51, x55_c, x56_c, x58, x59_c, x61, x62, x63_c, x64_c, x73, x74_c, x75_c, x76_c, x77_c, x79, x81_c, x82, x89, x90_c, x91_c, x93, x94_c, x96, x97_c, x98);
and (w6486, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x64, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6487, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47_c, x73_c, x76, x85, x89, x91_c, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6488, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6489, x0_c, x3, x4_c, x5, x6, x7, x8, x10_c, x11_c, x12_c, x13, x14, x17, x20_c, x22_c, x24_c, x27_c, x28_c, x29, x30_c, x31_c, x32, x38_c, x39, x40, x41, x42, x44, x45_c, x46_c, x50, x51_c, x55_c, x57, x59, x63, x70_c, x71, x72_c, x74_c, x75, x76, x77_c, x80_c, x82, x85, x86_c, x87, x88, x89, x90, x93, x94, x96, x97_c);
and (w6490, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x27, x57_c, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6491, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75, x83_c);
and (w6492, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6493, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x63, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6494, x0, x4_c, x12, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6495, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x95, x99);
and (w6496, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6497, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x85, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6498, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6499, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x52_c, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6500, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89_c, x93_c, x97_c);
and (w6501, x20, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6502, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6503, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6504, x0, x3, x6, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6505, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6506, x0, x4_c, x15_c, x22_c, x25_c, x29, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6507, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6508, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17_c, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6509, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21_c, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6510, x2_c, x7, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6511, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6512, x1, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6513, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x54, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6514, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6515, x2_c, x11, x29_c, x56_c, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6516, x0, x2, x3, x4_c, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6517, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6518, x2, x5, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6519, x0, x1_c, x3, x4, x5, x6, x8_c, x9, x10_c, x11, x12, x13_c, x15_c, x16, x17_c, x18, x19_c, x24, x25, x26, x27_c, x28, x29_c, x30_c, x32_c, x33, x34_c, x35_c, x36, x37, x38, x39_c, x40, x41_c, x42_c, x45_c, x46_c, x47, x49_c, x50, x51_c, x52, x53_c, x54, x55_c, x56_c, x58_c, x59, x60, x61, x62, x63, x64_c, x65, x67, x68, x69, x70, x71_c, x72_c, x73, x74_c, x76_c, x77_c, x78_c, x79_c, x80, x82, x83_c, x84_c, x85, x87, x88, x89_c, x90, x92, x93, x94_c, x96_c, x97, x98, x99);
and (w6520, x0, x2, x7_c, x8_c, x11_c, x15_c, x22_c, x25_c, x26, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6521, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87_c, x88, x89_c, x90_c, x91_c, x92, x93, x95, x96, x97_c, x98);
and (w6522, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6523, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6524, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60, x61_c, x63_c, x65, x72_c, x81, x84, x85, x95, x99);
and (w6525, x0, x1, x2, x3_c, x4, x6_c, x7_c, x8_c, x9, x10, x11_c, x12, x13, x14_c, x15, x18, x19, x20_c, x22_c, x23_c, x24_c, x25, x26, x28_c, x29, x32_c, x33, x34_c, x35_c, x36, x37, x38, x40, x42, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x51, x52, x53_c, x54_c, x55, x56_c, x57_c, x58, x59, x60_c, x61, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x71, x72, x74_c, x75_c, x76_c, x77, x79_c, x81, x82, x83_c, x84, x85, x86, x87, x88, x91, x92_c, x93, x96_c, x97_c, x98_c, x99);
and (w6526, x49, x94_c, x96_c, x97);
and (w6527, x0, x1, x2_c, x3_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6528, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x36_c, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6529, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6530, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x54, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6531, x1_c, x3_c, x4_c, x5_c, x6, x7, x8_c, x9, x10, x11_c, x13, x14, x16, x18, x19_c, x20, x21, x22_c, x23, x24, x25, x26_c, x27_c, x28, x30, x31_c, x32, x33_c, x35, x36_c, x37_c, x38_c, x40, x41_c, x42_c, x43, x44_c, x45_c, x46, x47_c, x48_c, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56_c, x57_c, x58_c, x59_c, x60, x62, x63_c, x64, x65, x66, x67, x69, x70, x71, x72, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x81, x82, x83_c, x84, x87_c, x88, x89_c, x91, x92_c, x94_c, x95, x96, x97, x98_c, x99_c);
and (w6532, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6533, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6534, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8, x9, x10, x11, x12, x13_c, x14_c, x15_c, x16, x17_c, x18, x19_c, x20_c, x21_c, x22, x23, x24, x25, x26, x27_c, x28_c, x29, x30, x31, x32_c, x33, x35_c, x36_c, x37, x38, x39_c, x40_c, x41_c, x42_c, x43, x44_c, x46, x47, x48, x49, x50_c, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70_c, x71_c, x72, x73_c, x74, x75, x76_c, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84, x85, x86_c, x87, x88_c, x89, x90_c, x91, x92_c, x93, x94, x95, x96_c, x97, x98);
and (w6535, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x45_c, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6536, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92, x93_c, x95_c, x96, x97, x98);
and (w6537, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x44_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6538, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6539, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89, x90_c, x94_c, x95, x96, x97_c);
and (w6540, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x65_c, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6541, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x75, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6542, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x63, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6543, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6544, x46, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6545, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x51_c, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6546, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x87, x88_c, x93_c, x97_c);
and (w6547, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42, x44_c, x57, x72, x73, x75_c, x76, x77, x78, x79, x80, x81_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6548, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6549, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6550, x0, x1, x2_c, x3, x4_c, x5_c, x6, x7_c, x8, x9_c, x10_c, x11_c, x12, x14_c, x15, x16_c, x17_c, x18_c, x19, x20_c, x21, x22, x24, x25, x26_c, x27_c, x28, x30, x31, x33_c, x34_c, x35_c, x37_c, x38, x39_c, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x49_c, x50_c, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61, x62, x66_c, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80_c, x81, x82_c, x83, x84, x85_c, x86_c, x87, x88_c, x89, x90_c, x92, x93_c, x94, x95, x97, x98_c, x99);
and (w6551, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6552, x0_c, x5, x23_c, x30_c, x31, x32, x35, x36, x37, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83_c, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6553, x0_c, x1, x2, x3, x4_c, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12, x13, x14, x15, x16, x17_c, x18, x19_c, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30_c, x31, x32, x33, x34, x35_c, x36_c, x37, x38, x39, x40_c, x41, x42, x43, x44_c, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58_c, x59_c, x60_c, x61, x62_c, x63, x64_c, x65, x66, x67_c, x68_c, x69_c, x70, x71_c, x72, x73, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81_c, x82_c, x83, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96_c, x97, x98, x99);
and (w6554, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x92_c, x95, x97_c);
and (w6555, x0, x6_c, x7_c, x9, x12_c, x14, x15, x17, x19, x20_c, x22_c, x23_c, x25, x26, x27, x28_c, x30_c, x34_c, x36, x37_c, x42, x43, x46, x47, x49_c, x53_c, x55, x56_c, x58_c, x61_c, x62_c, x64, x65_c, x67_c, x69_c, x74_c, x76, x77, x78_c, x81, x82, x83_c, x84_c, x86_c, x87_c, x89_c, x91_c, x92_c, x94, x95, x96_c, x98_c, x99_c);
and (w6556, x11_c, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6557, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w6558, x3_c, x8_c, x14, x23_c, x24, x29, x31, x36, x47_c, x53_c, x58, x69, x74, x78_c, x80_c, x86, x87_c, x88, x89, x90, x98_c);
and (w6559, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x42_c, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6560, x2_c, x6_c, x8, x10_c, x11_c, x14_c, x17, x18_c, x22_c, x24, x25_c, x31, x33_c, x38_c, x41, x47, x49_c, x50_c, x52, x58, x60, x62_c, x65_c, x71_c, x74, x75_c, x77, x78_c, x81, x84, x89_c, x95_c, x96);
and (w6561, x8, x21_c, x25_c, x26, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6562, x0, x3, x4, x5, x6_c, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6563, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x56, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6564, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6565, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x70_c, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6566, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x80_c, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6567, x9_c, x12, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6568, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x46, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x89, x93, x97_c, x98_c, x99_c);
and (w6569, x0, x7, x8_c, x10, x15_c, x26, x35, x36_c, x38, x40_c, x41, x43, x52, x59_c, x61, x63_c, x65_c, x66, x68_c, x70, x71, x73, x76, x78_c, x84, x85, x88_c, x93, x99);
and (w6570, x0, x1, x2, x3_c, x4, x6, x9, x10_c, x11_c, x12_c, x13_c, x14_c, x17, x19, x20_c, x21_c, x22, x23, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x35, x36, x37_c, x38, x39, x40_c, x41_c, x43, x44_c, x45_c, x46_c, x47, x48_c, x49, x51_c, x52, x53, x54_c, x55_c, x58, x60_c, x61, x62, x64, x65_c, x67, x68_c, x69_c, x70_c, x71, x72, x74_c, x76_c, x77_c, x78_c, x79, x80_c, x81_c, x82, x83, x84, x85, x86_c, x87, x88_c, x89_c, x91, x92, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6571, x0, x3, x10, x13, x14, x15, x16_c, x22, x32_c, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6572, x0, x1_c, x2, x3, x5_c, x6_c, x7, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6573, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6574, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6575, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6576, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70_c, x73_c, x76, x85, x86, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6577, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35_c, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6578, x0_c, x1, x2, x3_c, x4_c, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6579, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6580, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6581, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x76, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6582, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6583, x12_c, x38, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60_c, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6584, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6585, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6586, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6587, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6588, x0_c, x1_c, x2, x3_c, x5_c, x6_c, x7, x11_c, x12_c, x13, x15, x17_c, x18_c, x19_c, x20_c, x21_c, x25_c, x28_c, x33_c, x35, x37, x38_c, x39_c, x42_c, x44, x50, x51_c, x52_c, x53, x54_c, x56_c, x57, x58_c, x59, x60_c, x63, x64_c, x65, x66, x67_c, x68, x74_c, x76_c, x77, x78, x79_c, x82, x83, x84_c, x85, x88, x89, x90, x95_c, x96, x98_c, x99);
and (w6589, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44_c, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6590, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6591, x49, x84, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6592, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x50, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6593, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x37, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6594, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6595, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36, x83_c, x89_c, x93_c, x95_c, x96_c, x97_c);
and (w6596, x0, x1, x2, x3, x4_c, x6_c, x7, x10, x11_c, x13, x14_c, x15, x16, x17_c, x18, x20_c, x21_c, x22_c, x23_c, x25, x26, x27, x29_c, x30_c, x31, x35_c, x36, x37_c, x39, x40, x41, x42, x43_c, x45, x46_c, x47_c, x49_c, x52_c, x54, x58_c, x59, x60, x61, x62, x64_c, x65_c, x68, x69_c, x70_c, x71, x72, x73, x74, x76_c, x77_c, x78_c, x82, x83, x84_c, x86_c, x87_c, x88_c, x89, x90_c, x91, x92, x96_c, x97_c, x98, x99);
and (w6597, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x77, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6598, x0, x1_c, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w6599, x0, x1, x2_c, x3, x4_c, x5, x6, x7_c, x8_c, x10_c, x12_c, x14_c, x17, x18_c, x20_c, x21_c, x22_c, x24, x27, x28, x29_c, x31_c, x32_c, x35, x36, x37, x38_c, x39, x41_c, x42, x43_c, x44_c, x45, x47, x49_c, x50_c, x51_c, x53, x54, x56, x57, x58_c, x59, x60_c, x62_c, x65_c, x66, x68, x69_c, x70, x71_c, x72, x73, x74_c, x76, x77_c, x81_c, x83, x84, x85_c, x86, x87_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98_c);
and (w6600, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6601, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6602, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84_c, x87, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6603, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6604, x0_c, x2_c, x3_c, x5_c, x6_c, x8, x9_c, x10, x11_c, x12, x13_c, x14, x15_c, x16_c, x18, x19, x20_c, x21_c, x22, x23, x24, x25, x26_c, x27_c, x28_c, x29_c, x30, x31_c, x32, x33_c, x34, x35, x36, x37, x38_c, x39, x41_c, x42_c, x43, x44, x45_c, x47, x48_c, x49, x50_c, x51, x53, x54_c, x55_c, x57_c, x58, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66, x67, x69_c, x70_c, x71, x73_c, x74, x75, x76, x79, x80_c, x82_c, x83, x84, x85, x88_c, x89_c, x90, x91_c, x93, x95_c, x96_c, x97, x98, x99_c);
and (w6605, x0, x1_c, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6606, x40_c, x56, x92_c);
and (w6607, x0, x3, x10, x13, x14, x15, x16_c, x18_c, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6608, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7, x8, x9_c, x10, x11_c, x12_c, x13, x14, x16_c, x17_c, x18, x19, x20_c, x21, x22, x23, x24_c, x26, x27_c, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x41_c, x42, x43, x44, x45, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55_c, x56, x57_c, x59_c, x60_c, x61, x62, x63_c, x64_c, x65, x66, x67_c, x68, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x76_c, x77_c, x78, x79_c, x80, x81_c, x82, x83, x84_c, x86, x87, x88, x89, x90, x91, x92_c, x93_c, x94, x95_c, x96, x97, x98_c);
and (w6609, x0_c, x1_c, x4_c, x5, x6_c, x8, x10_c, x12_c, x13_c, x15, x16_c, x18, x22_c, x23, x25, x26_c, x27_c, x32_c, x36_c, x37, x38, x39, x40_c, x41_c, x43_c, x44, x45, x46, x47, x48_c, x51, x53, x54_c, x55_c, x57_c, x58_c, x60_c, x63, x65_c, x69_c, x70, x71_c, x72, x76_c, x77_c, x78_c, x80, x81_c, x82, x83_c, x85, x87_c, x96_c, x97_c);
and (w6610, x0, x1, x2_c, x3, x4, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x67_c, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6611, x5, x6, x7_c, x10, x11_c, x13, x20_c, x24, x29, x32_c, x37_c, x39_c, x40, x41_c, x44, x45, x46_c, x47, x52_c, x59_c, x60_c, x61_c, x63_c, x66_c, x67, x70, x72, x79, x81_c, x84_c, x85, x88, x89, x91, x96, x99_c);
and (w6612, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27, x83_c);
and (w6613, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x84_c, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6614, x0_c, x4_c, x5_c, x6_c, x8_c, x11, x12_c, x15_c, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x49, x64, x71, x72_c, x79, x85, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6615, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w6616, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w6617, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x86, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6618, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6619, x84_c, x90_c);
and (w6620, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x93, x95_c, x96, x98, x99);
and (w6621, x0_c, x3_c, x4_c, x10_c, x11, x13_c, x16, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6622, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x50, x51, x52_c, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6623, x6, x17_c, x20_c, x24_c, x25_c, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6624, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x58_c, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w6625, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92, x93, x94_c, x96_c, x97_c, x98);
and (w6626, x0_c, x1_c, x2, x3, x4, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13, x14_c, x15_c, x17_c, x18, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34_c, x35, x36, x37_c, x38, x39, x40, x42, x43, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x52, x53, x54, x55_c, x56_c, x57_c, x58, x59, x60, x62_c, x63, x64_c, x65, x66, x67, x69_c, x70_c, x71_c, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x82_c, x83, x84, x85_c, x86_c, x87, x88, x89_c, x91, x92, x93_c, x95_c, x96_c, x97, x98, x99);
and (w6627, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x45_c, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x87_c, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6628, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55_c, x83_c);
and (w6629, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x93, x97_c);
and (w6630, x0, x1, x3, x4_c, x5, x6, x7, x8_c, x9_c, x11_c, x12_c, x13, x14, x15, x18_c, x19_c, x20_c, x22, x23, x24, x25, x27, x28, x29_c, x30, x31, x32_c, x33_c, x34, x35_c, x38_c, x39, x40, x41, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49, x50_c, x51, x52, x53_c, x55_c, x56_c, x57, x58_c, x59_c, x60, x61_c, x62_c, x63, x65_c, x66, x67_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x79, x80, x81, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89, x90, x91, x92_c, x94_c, x95, x96_c, x97, x99_c);
and (w6631, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x44_c, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x82_c, x88_c, x93_c, x95_c);
and (w6632, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x83, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6633, x5_c, x9, x27, x61_c, x70_c, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6634, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x69_c, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x93, x95_c, x96, x98, x99);
and (w6635, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8, x9, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6636, x13_c, x49, x64, x72_c, x73, x75, x81_c, x87, x90, x93_c, x97_c);
and (w6637, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w6638, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89, x93_c, x97_c);
and (w6639, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6640, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6641, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x28, x29, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6642, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6643, x11, x12_c, x15, x16, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6644, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6645, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x45, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6646, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x22, x23_c, x24, x25_c, x26_c, x27, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6647, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6648, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6649, x0, x4_c, x6_c, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6650, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6651, x2, x3_c, x4, x6, x9, x10_c, x11_c, x12, x18, x19_c, x21_c, x22, x23, x25, x26, x30_c, x34_c, x35, x39_c, x40_c, x42_c, x43_c, x45, x47_c, x54_c, x58_c, x59, x63_c, x66_c, x67_c, x69_c, x70, x72, x78_c, x81, x83, x84_c, x85_c, x86_c, x94, x95_c, x98_c);
and (w6652, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6653, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x57, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6654, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88, x90_c, x91, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6655, x5_c, x8_c, x9, x11, x12_c, x13, x14_c, x15_c, x16_c, x19_c, x21_c, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37, x38, x40, x45, x46_c, x47, x49, x50, x51_c, x55_c, x56, x57_c, x58, x59_c, x60, x62, x64, x65_c, x66, x68_c, x69_c, x70_c, x71, x72_c, x74_c, x76_c, x77, x78_c, x81, x85, x87_c, x88, x90, x91, x93, x94_c, x95, x97_c, x98_c, x99_c);
and (w6656, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92_c, x93_c, x95_c, x96, x98, x99);
and (w6657, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6658, x1, x2, x4, x9, x11, x12, x17, x21, x22_c, x23, x24, x26, x34, x35_c, x36, x37_c, x38_c, x39, x40, x41_c, x43_c, x44, x46_c, x49, x51, x54_c, x65, x66_c, x68_c, x72_c, x80, x85, x91_c, x93_c, x94, x95, x96_c, x98);
and (w6659, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x95, x96, x97, x99_c);
and (w6660, x2_c, x11, x29_c, x44, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6661, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x26_c, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6662, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6663, x1, x4, x6, x8_c, x9_c, x10, x11, x13_c, x14, x15, x16, x18, x19_c, x20_c, x21_c, x22, x24, x25_c, x26, x27, x30, x31_c, x32_c, x36_c, x39_c, x40_c, x41_c, x42_c, x43, x46_c, x48, x49_c, x50_c, x52_c, x54, x55, x57_c, x58, x59, x63, x64_c, x67_c, x70, x71_c, x72_c, x74, x77, x79_c, x81, x82_c, x83, x84_c, x87_c, x88, x89_c, x91, x93_c, x94, x95, x98, x99_c);
and (w6664, x1, x11, x12_c, x15, x17_c, x22, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6665, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x51_c, x52_c, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6666, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6667, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6668, x2, x3_c, x4_c, x6_c, x7_c, x8_c, x10, x14, x15, x16, x18, x20, x21, x22_c, x25_c, x29, x31_c, x32_c, x33, x34_c, x35_c, x39_c, x41_c, x42_c, x44, x45_c, x46, x47, x48, x49, x50_c, x51_c, x52_c, x54, x55_c, x56_c, x58, x59, x60, x61_c, x62_c, x64_c, x67_c, x69_c, x73_c, x76_c, x78_c, x84, x86, x90_c, x91_c, x95, x96, x98_c);
and (w6669, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6670, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90);
and (w6671, x0, x1, x3, x10, x13, x14, x15, x16_c, x22, x33_c, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6672, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6673, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98_c);
and (w6674, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44_c, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6675, x0, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x80_c, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6676, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x83, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6677, x0_c, x1_c, x3, x4_c, x5, x7, x8_c, x9, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6678, x13_c, x49, x64, x71, x72_c, x79, x97);
and (w6679, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x69, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6680, x0, x1, x2_c, x3, x4, x5_c, x6, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32, x83_c);
and (w6681, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x62_c, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6682, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49, x73_c, x76, x85, x89, x93, x97_c);
and (w6683, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6684, x0, x2_c, x5_c, x12, x13, x14_c, x16, x24, x25_c, x26, x30, x33_c, x34_c, x40_c, x43, x44_c, x45, x46, x53_c, x58, x59_c, x61, x63_c, x68, x69, x75_c, x77, x78, x79_c, x80, x81, x83_c, x85, x87, x89, x90, x92, x93_c, x94_c, x98);
and (w6685, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26_c, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96, x97_c);
and (w6686, x5_c, x9, x27, x61_c, x76, x88_c, x95_c, x97_c);
and (w6687, x4_c, x10, x15_c, x16_c, x21_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6688, x6, x10, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w6689, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91, x92, x93_c, x94, x95_c, x96, x99_c);
and (w6690, x12_c, x32, x68_c, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6691, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x44, x47_c, x49_c, x56, x60, x61_c, x63_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6692, x49, x72, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95, x97_c);
and (w6693, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95_c, x97_c);
and (w6694, x0_c, x5, x23_c, x30_c, x31, x32, x36_c, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6695, x4_c, x10, x15_c, x22_c, x24_c, x25_c, x32_c, x34_c, x35, x41, x42_c, x44_c, x47_c, x49_c, x56, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6696, x0_c, x2, x6, x9_c, x15, x17, x21_c, x22, x24, x26_c, x27, x29, x30_c, x32, x38_c, x40_c, x41, x44_c, x45, x47, x48, x49_c, x50, x52_c, x53, x54_c, x58_c, x60, x61_c, x64, x67, x69, x71_c, x72, x73, x74_c, x77, x78, x79_c, x87, x88_c, x89, x90, x91_c, x93, x95, x96_c);
and (w6697, x2_c, x8_c, x15_c, x26, x35, x36, x51, x54_c, x69_c, x70, x71, x77, x79, x82_c, x84_c, x93_c, x94, x95, x96_c, x98);
and (w6698, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73);
and (w6699, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39_c, x71_c);
and (w6700, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6701, x8, x9_c, x14_c, x15_c, x21_c, x25_c, x31_c, x36_c, x39_c, x42_c, x46, x60, x61, x62, x67, x69_c, x73_c, x74_c, x75_c, x76, x77, x79_c, x83, x84, x85_c, x86_c, x88, x89_c, x90_c, x93_c, x95, x96, x97);
and (w6702, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57_c, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6703, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x18, x19_c, x21, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6704, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6705, x1_c, x10, x15_c, x17, x19_c, x24_c, x27_c, x32_c, x46, x49, x70_c, x75_c, x81, x83_c, x90_c, x98_c);
and (w6706, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x47, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6707, x27_c, x28, x29_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6708, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w6709, x0, x6_c, x12, x13_c, x15_c, x17_c, x18_c, x19_c, x20, x22_c, x23, x25_c, x29_c, x30, x32, x35, x40_c, x41_c, x45_c, x46, x47, x49_c, x50, x52, x56, x58_c, x60_c, x62, x64, x65, x66, x68, x71_c, x72_c, x76, x77, x78, x79_c, x88_c, x89_c, x90_c, x91, x92, x93_c, x97_c, x99);
and (w6710, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x32_c, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w6711, x9_c, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6712, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10, x13, x16_c, x17, x18, x26, x27, x28_c, x33, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51_c, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6713, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6714, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6715, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x93_c, x95_c, x97, x98_c, x99_c);
and (w6716, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6717, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6718, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6719, x12_c, x32, x91, x95_c, x96, x97_c, x98, x99);
and (w6720, x0_c, x4_c, x5, x13_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6721, x12_c, x25, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6722, x10_c, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6723, x1, x5, x9_c, x12, x13, x15_c, x17, x22_c, x25_c, x31_c, x40_c, x47_c, x48, x51, x61_c, x62_c, x65, x66, x72_c, x74_c, x76_c, x80, x84, x85_c);
and (w6724, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x17, x18, x20, x21, x23_c, x25, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6725, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6726, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x77, x78_c, x79_c, x81_c, x82, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6727, x0_c, x4_c, x5_c, x6, x13_c, x49, x64, x71, x72_c, x79, x90_c, x93_c, x97_c);
and (w6728, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6729, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x66, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6730, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72, x73_c, x76, x85, x89, x93, x97_c);
and (w6731, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x47_c, x49_c, x56, x60, x61_c, x65_c, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6732, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6733, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x21, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6734, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80_c, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6735, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6736, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81_c, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w6737, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x61_c, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w6738, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16_c, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x81_c, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6739, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89, x93, x97_c);
and (w6740, x12_c, x32, x35, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w6741, x0_c, x1, x2_c, x3, x4_c, x5, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6742, x49, x76, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w6743, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6744, x2, x6_c, x7_c, x8, x10, x12_c, x13, x14_c, x15, x17, x19_c, x20_c, x22, x23_c, x24, x25, x29, x30, x34, x36, x40_c, x42_c, x50_c, x51, x52, x55_c, x56_c, x57, x58, x59_c, x60_c, x61, x62_c, x65, x66, x67, x69, x75, x79, x80_c, x81_c, x82_c, x89, x91, x92, x95_c, x96, x97);
and (w6745, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x82_c, x83_c, x85_c, x86_c, x87_c, x88, x90, x93_c, x95_c, x96, x98, x99);
and (w6746, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38, x39, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x99_c);
and (w6747, x0, x2_c, x5, x10, x16, x21_c, x31, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w6748, x9_c, x10_c, x16_c, x25_c, x44_c, x50, x57, x63_c, x64_c, x65, x68_c, x70, x83_c, x89, x92_c);
and (w6749, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23, x25_c, x27, x31, x33, x34_c, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x58, x59_c, x60, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w6750, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w6751, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47_c, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w6752, x0, x1_c, x5_c, x9, x27, x53_c, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6753, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89, x90_c, x92, x93_c, x94_c, x95, x96_c, x97, x98, x99_c);
and (w6754, x7, x9, x10_c, x12, x14_c, x18_c, x19_c, x22, x23, x24, x26, x27, x34, x40, x46_c, x48_c, x53, x55, x57_c, x62, x63_c, x65, x70_c, x71, x72, x73, x74_c, x79, x80, x84, x86, x87_c, x89, x90, x92, x98_c, x99);
and (w6755, x8, x21_c, x25_c, x27_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x82, x84_c, x86_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w6756, x1_c, x2, x4, x5, x6_c, x8_c, x9, x11_c, x13, x14_c, x16_c, x19, x20_c, x21, x22_c, x23_c, x24, x25, x26_c, x27_c, x29_c, x30_c, x31, x33, x34_c, x35, x36, x40, x41_c, x42_c, x43, x44, x45, x46, x47, x48, x50_c, x52_c, x53, x55_c, x57_c, x59, x61_c, x62_c, x63_c, x65_c, x66, x67, x70, x71, x72, x73_c, x74, x75, x76_c, x77_c, x79, x82, x83_c, x85_c, x90, x91, x92, x94_c, x95_c, x96, x97_c, x98_c, x99);
and (w6757, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x30, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75_c, x86, x89_c, x90_c, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
xor (o, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757);
endmodule
