module top(x0, x1, x2, x3, x4, x5, x6, x7,  o);
input x0, x1, x2, x3, x4, x5, x6, x7;
output o;
wire x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9;
assign x0_c = ~x0;
assign x1_c = ~x1;
assign x2_c = ~x2;
assign x3_c = ~x3;
assign x4_c = ~x4;
assign x5_c = ~x5;
assign x6_c = ~x6;
assign x7_c = ~x7;
and (w0, x1_c, x2, x3_c, x4, x5_c, x6_c, x7);
and (w1, x0, x1_c, x2, x3, x4_c, x5_c, x6, x7);
and (w2, x4_c, x5_c, x6_c);
and (w3, x1, x3, x5, x7);
and (w4, x0, x1_c, x2, x3, x4, x5_c, x6_c);
and (w5, x1_c, x2, x3, x5, x6_c, x7_c);
and (w6, x6, x7);
and (w7, x0_c, x2, x4, x7_c);
and (w8, x0, x1_c, x2_c);
assign w9 = x5_c;
xor (o, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9);
endmodule
