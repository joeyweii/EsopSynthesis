module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,  o);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
output o;
wire x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70;
assign x0_c = ~x0;
assign x1_c = ~x1;
assign x2_c = ~x2;
assign x3_c = ~x3;
assign x4_c = ~x4;
assign x5_c = ~x5;
assign x6_c = ~x6;
assign x7_c = ~x7;
assign x8_c = ~x8;
assign x9_c = ~x9;
and (w0, x6, x8);
and (w1, x0, x2_c, x4_c, x5_c, x6, x7, x8, x9_c);
and (w2, x1_c, x8, x9_c);
and (w3, x2, x3, x4_c, x5_c, x6, x7_c, x8, x9_c);
and (w4, x3, x4, x9);
and (w5, x0, x4_c);
and (w6, x0, x1_c, x2, x3_c, x5, x7, x8_c);
and (w7, x0_c, x1);
and (w8, x0_c, x3, x4, x6, x9_c);
and (w9, x0, x1_c, x2_c, x3_c, x7);
assign w10 = x7;
and (w11, x1_c, x2, x6_c, x7, x8_c);
and (w12, x0, x2_c, x7);
and (w13, x1_c, x2, x4, x8_c, x9);
and (w14, x2_c, x5, x6, x7_c, x8, x9);
and (w15, x4_c, x7);
and (w16, x0, x1_c, x2, x3_c, x4, x5_c, x6_c, x7, x8_c, x9);
and (w17, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7, x8_c, x9);
and (w18, x0, x2, x3, x4, x5, x6, x7_c, x8);
and (w19, x0_c, x1_c, x2, x4_c, x5_c, x6_c, x7, x8_c, x9);
and (w20, x1_c, x3, x4_c, x5_c, x8_c, x9_c);
and (w21, x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x8);
and (w22, x0, x1, x2_c, x3, x4_c, x5_c, x6, x7, x8, x9_c);
and (w23, x0, x2_c, x3_c, x4, x5, x7_c);
and (w24, x0, x1, x2_c, x7_c, x9_c);
and (w25, x0, x1_c, x2_c, x3, x5_c, x6_c, x7, x8_c, x9_c);
and (w26, x3_c, x4, x6, x7_c);
and (w27, x0_c, x1_c, x2, x4_c, x5, x6_c, x7, x8, x9_c);
and (w28, x1, x2_c, x4, x6, x7, x8_c);
and (w29, x0_c, x3_c, x4_c, x5, x6_c, x7_c, x9_c);
and (w30, x1_c, x2_c, x4, x5_c, x8_c, x9);
and (w31, x0_c, x1_c, x2, x3_c, x4, x5, x6, x8, x9);
and (w32, x0_c, x1, x3_c, x4_c, x5, x6_c, x7, x8_c, x9_c);
and (w33, x1_c, x2_c, x4, x6, x7_c, x8);
and (w34, x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c);
and (w35, x0_c, x3, x6, x8_c, x9);
and (w36, x0, x1_c, x2, x3, x4, x5_c, x6, x7_c, x8_c, x9_c);
and (w37, x4_c, x8);
and (w38, x2, x6_c);
and (w39, x0, x1_c, x2_c, x3, x4_c, x5_c, x6_c, x7_c, x9);
and (w40, x3, x4_c, x8_c);
and (w41, x0, x2, x3, x5, x6, x7, x8, x9);
and (w42, x0, x1_c, x2, x3_c, x4_c, x5, x6_c, x7, x8_c, x9);
and (w43, x0_c, x4, x6_c, x8_c, x9);
and (w44, x1_c, x2, x4, x5, x9_c);
and (w45, x0_c, x2, x4, x6_c);
and (w46, x0, x1_c, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9);
and (w47, x2_c, x7_c, x9);
and (w48, x1_c, x3_c, x4_c, x5, x6_c, x7, x9_c);
and (w49, x0_c, x1_c, x3, x4_c, x8, x9_c);
and (w50, x0, x2_c, x4_c, x8_c, x9);
and (w51, x2, x3_c, x5_c, x6, x7, x8, x9);
and (w52, x2, x3_c, x6_c, x7, x8_c, x9);
and (w53, x0, x1, x2_c, x4, x9);
and (w54, x5_c, x6_c);
and (w55, x0, x3, x4_c, x7_c);
and (w56, x1_c, x3_c, x4_c, x7, x8, x9_c);
assign w57 = x1;
and (w58, x3_c, x6, x8_c);
and (w59, x0, x1, x2, x3, x4_c, x5, x6_c, x7, x8_c, x9_c);
and (w60, x1, x2_c, x3, x4_c, x5_c, x6_c, x7, x8, x9_c);
and (w61, x1_c, x2_c, x3, x4_c, x5_c, x9);
and (w62, x1, x2_c, x4, x6_c);
and (w63, x1, x3, x5_c, x7);
and (w64, x0_c, x1_c, x2_c, x3_c, x4_c, x6);
and (w65, x1_c, x2, x4_c, x6, x7);
and (w66, x0, x1_c, x3_c);
and (w67, x0, x1, x2, x3_c, x4_c, x5, x6_c, x7, x8_c, x9_c);
and (w68, x0, x1_c, x2_c, x3_c, x4_c, x6);
assign w69 = x0_c;
and (w70, x0, x1_c, x2_c, x3, x4, x7_c, x8_c, x9_c);
xor (o, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70);
endmodule
