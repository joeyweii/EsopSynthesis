module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,  o);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
output o;
wire x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19;
assign x0_c = ~x0;
assign x1_c = ~x1;
assign x2_c = ~x2;
assign x3_c = ~x3;
assign x4_c = ~x4;
assign x5_c = ~x5;
assign x6_c = ~x6;
assign x7_c = ~x7;
assign x8_c = ~x8;
assign x9_c = ~x9;
assign w0 = x9;
and (w1, x3_c, x5, x6, x7_c, x8, x9_c);
and (w2, x3_c, x4_c);
and (w3, x1_c, x3_c, x4_c, x5, x6, x8_c, x9_c);
and (w4, x1, x3, x4_c, x6, x7, x8_c, x9);
and (w5, x0, x4_c, x6, x9_c);
and (w6, x1_c, x2_c, x3, x4_c, x5_c, x6_c, x7_c, x8_c, x9);
and (w7, x0_c, x1_c, x2, x3_c, x4_c, x5_c, x6_c, x8_c);
and (w8, x0_c, x1, x2_c, x7, x9);
and (w9, x0_c, x3_c, x4_c, x5, x6, x7_c, x8_c, x9);
and (w10, x1_c, x2);
and (w11, x3, x5_c, x6_c, x9);
and (w12, x2_c, x4_c, x5_c, x9);
and (w13, x0, x1_c, x6_c, x7);
and (w14, x0, x1, x3, x4, x6_c, x7, x8_c);
and (w15, x3, x4_c, x5_c, x8);
and (w16, x0, x1_c, x2_c, x3, x4_c, x5, x6_c, x7, x8_c, x9);
and (w17, x1_c, x3, x4, x9_c);
and (w18, x0_c, x1_c, x2, x3, x4, x5, x6_c, x7_c, x9_c);
and (w19, x0_c, x1_c, x2_c, x3_c, x4, x5, x6_c, x7, x8, x9);
xor (o, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19);
endmodule
