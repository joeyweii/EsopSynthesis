module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99,  o);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99;
output o;
wire x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31_c, x32_c, x33_c, x34_c, x35_c, x36_c, x37_c, x38_c, x39_c, x40_c, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98_c, x99_c;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999;
assign x0_c = ~x0;
assign x1_c = ~x1;
assign x2_c = ~x2;
assign x3_c = ~x3;
assign x4_c = ~x4;
assign x5_c = ~x5;
assign x6_c = ~x6;
assign x7_c = ~x7;
assign x8_c = ~x8;
assign x9_c = ~x9;
assign x10_c = ~x10;
assign x11_c = ~x11;
assign x12_c = ~x12;
assign x13_c = ~x13;
assign x14_c = ~x14;
assign x15_c = ~x15;
assign x16_c = ~x16;
assign x17_c = ~x17;
assign x18_c = ~x18;
assign x19_c = ~x19;
assign x20_c = ~x20;
assign x21_c = ~x21;
assign x22_c = ~x22;
assign x23_c = ~x23;
assign x24_c = ~x24;
assign x25_c = ~x25;
assign x26_c = ~x26;
assign x27_c = ~x27;
assign x28_c = ~x28;
assign x29_c = ~x29;
assign x30_c = ~x30;
assign x31_c = ~x31;
assign x32_c = ~x32;
assign x33_c = ~x33;
assign x34_c = ~x34;
assign x35_c = ~x35;
assign x36_c = ~x36;
assign x37_c = ~x37;
assign x38_c = ~x38;
assign x39_c = ~x39;
assign x40_c = ~x40;
assign x41_c = ~x41;
assign x42_c = ~x42;
assign x43_c = ~x43;
assign x44_c = ~x44;
assign x45_c = ~x45;
assign x46_c = ~x46;
assign x47_c = ~x47;
assign x48_c = ~x48;
assign x49_c = ~x49;
assign x50_c = ~x50;
assign x51_c = ~x51;
assign x52_c = ~x52;
assign x53_c = ~x53;
assign x54_c = ~x54;
assign x55_c = ~x55;
assign x56_c = ~x56;
assign x57_c = ~x57;
assign x58_c = ~x58;
assign x59_c = ~x59;
assign x60_c = ~x60;
assign x61_c = ~x61;
assign x62_c = ~x62;
assign x63_c = ~x63;
assign x64_c = ~x64;
assign x65_c = ~x65;
assign x66_c = ~x66;
assign x67_c = ~x67;
assign x68_c = ~x68;
assign x69_c = ~x69;
assign x70_c = ~x70;
assign x71_c = ~x71;
assign x72_c = ~x72;
assign x73_c = ~x73;
assign x74_c = ~x74;
assign x75_c = ~x75;
assign x76_c = ~x76;
assign x77_c = ~x77;
assign x78_c = ~x78;
assign x79_c = ~x79;
assign x80_c = ~x80;
assign x81_c = ~x81;
assign x82_c = ~x82;
assign x83_c = ~x83;
assign x84_c = ~x84;
assign x85_c = ~x85;
assign x86_c = ~x86;
assign x87_c = ~x87;
assign x88_c = ~x88;
assign x89_c = ~x89;
assign x90_c = ~x90;
assign x91_c = ~x91;
assign x92_c = ~x92;
assign x93_c = ~x93;
assign x94_c = ~x94;
assign x95_c = ~x95;
assign x96_c = ~x96;
assign x97_c = ~x97;
assign x98_c = ~x98;
assign x99_c = ~x99;
and (w0, x0, x6, x14_c, x16, x18, x19_c, x20, x22_c, x24, x25_c, x32_c, x41_c, x43_c, x46_c, x48_c, x49, x51, x55_c, x59_c, x61_c, x66, x68, x75_c, x76, x79, x80_c, x84, x85, x88, x91_c, x93);
and (w1, x4_c, x5_c, x7_c, x8, x9_c, x10_c, x11_c, x14_c, x15_c, x16, x17, x21_c, x22_c, x24, x25_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x35, x36_c, x37, x38, x41, x45_c, x46_c, x47_c, x52, x53, x54_c, x56_c, x60, x61, x64_c, x67, x68, x69, x71_c, x75_c, x76, x78, x79_c, x81_c, x84_c, x87, x88, x89, x91_c, x92_c, x94, x95_c, x97, x99);
and (w2, x2, x3_c, x4, x6_c, x8, x10, x12_c, x13_c, x16, x19, x21, x22_c, x23_c, x25, x26_c, x28, x29_c, x30, x31_c, x34, x35, x36_c, x39, x41, x42_c, x43_c, x44_c, x45_c, x50, x51, x52, x55, x59_c, x61_c, x62_c, x64, x65_c, x67_c, x68_c, x70_c, x71, x72, x73_c, x74, x75, x76, x77_c, x79, x80_c, x81, x82_c, x83, x86, x87, x88, x89, x91, x92, x93, x94_c, x97, x99);
and (w3, x17, x30, x38, x41_c, x72, x83_c, x91);
and (w4, x1_c, x2, x4, x5, x6_c, x9_c, x10, x11, x12_c, x14_c, x17, x18_c, x20_c, x21, x22_c, x25, x26_c, x28, x30, x31_c, x32, x34_c, x35_c, x37, x38, x42_c, x46, x47, x48_c, x52_c, x54_c, x57, x59_c, x60, x64_c, x66, x67, x68, x70_c, x73, x75_c, x77, x84_c, x85, x86, x87_c, x88, x90_c, x91, x94, x95_c, x98_c, x99_c);
and (w5, x2, x3, x7_c, x14_c, x17_c, x22, x23, x24, x26, x27, x31, x33, x35_c, x38, x39_c, x41, x42_c, x46, x48_c, x49, x54_c, x56, x57, x58_c, x62_c, x65_c, x71, x72, x79, x82_c, x84_c, x89_c, x90_c, x91_c, x97);
and (w6, x1, x5, x9_c, x12, x13, x15_c, x17, x22_c, x25_c, x31_c, x40_c, x47_c, x48, x51, x61_c, x62_c, x65, x66, x72_c, x74_c, x76_c, x80, x84, x85_c);
and (w7, x2_c, x3_c, x5_c, x6_c, x7_c, x8_c, x10, x11, x12, x15, x16, x17, x22_c, x25, x28_c, x29_c, x31, x33, x38_c, x39, x42_c, x45, x46_c, x47, x50_c, x51, x54_c, x55, x56, x58, x60, x61, x64, x65, x66, x70_c, x71_c, x72_c, x75_c, x78, x81, x82_c, x84_c, x85, x88, x89_c, x92_c, x93, x95_c, x96_c, x97, x98, x99);
and (w8, x3_c, x10_c, x14_c, x21_c, x29, x34_c, x41_c, x43, x81, x84_c, x86, x99_c);
and (w9, x0_c, x1_c, x3, x4_c, x5_c, x6_c, x7_c, x8, x9_c, x11, x12_c, x13_c, x14, x15_c, x18, x20, x21_c, x22, x24, x26, x27, x30, x37_c, x38, x39, x40_c, x41, x42_c, x43, x46, x47, x50_c, x52_c, x55, x58, x61_c, x63_c, x64_c, x67, x69, x71, x74, x76, x78_c, x80_c, x81_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91, x92, x94_c, x96, x98, x99_c);
and (w10, x8_c, x12_c, x14, x15, x18_c, x19, x23_c, x24_c, x26, x30, x32, x35, x36_c, x41_c, x47_c, x56_c, x76_c, x77_c, x78_c, x82, x90, x91_c, x98, x99);
and (w11, x2_c, x12, x16_c, x17_c, x18_c, x25, x29, x34_c, x40_c, x41_c, x44, x46_c, x50_c, x51_c, x53_c, x56, x58_c, x59, x60, x61_c, x65_c, x66_c, x71_c, x80_c, x82_c, x83, x84, x87, x91_c, x93_c, x95_c, x96_c);
and (w12, x1_c, x24_c, x31_c, x39_c, x47, x55_c, x58, x63_c, x73_c, x78_c, x80_c, x85, x89_c, x92_c, x94);
and (w13, x0, x37, x49, x85_c);
and (w14, x3, x13, x24, x27_c, x29, x31_c, x33_c, x35_c, x38_c, x41, x42, x53, x54_c, x57_c, x59, x61_c, x67, x68, x74, x75_c, x77_c, x78, x81, x85_c, x86, x90, x99);
and (w15, x1_c, x7, x8, x12, x15, x17, x20_c, x23, x24_c, x27_c, x32_c, x35_c, x36_c, x39, x40_c, x43, x49, x51_c, x53, x55_c, x59_c, x63_c, x65, x69_c, x70, x72, x76_c, x82_c, x83_c, x85_c, x87, x89_c, x92, x93, x96_c, x97);
and (w16, x1, x2_c, x5_c, x6_c, x9_c, x14_c, x17, x18_c, x19, x24, x27_c, x31, x37_c, x40, x41, x46, x49, x51, x61, x68, x90_c, x96_c);
and (w17, x0, x1, x2_c, x4_c, x5, x6, x7_c, x9_c, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x18, x19, x20, x22_c, x23, x25, x27, x28, x29_c, x30_c, x31, x32, x33_c, x34_c, x35_c, x37, x39, x40, x41_c, x42_c, x43, x44_c, x45_c, x46, x47_c, x48_c, x50, x51_c, x52, x53, x54, x55_c, x56, x57_c, x58_c, x59, x60, x61_c, x62_c, x64, x65_c, x66_c, x70, x71_c, x73, x75_c, x77_c, x78_c, x79, x81, x82_c, x83_c, x89, x90_c, x91_c, x93, x95, x96_c, x97, x99);
and (w18, x0, x1_c, x3_c, x4_c, x6, x7, x8_c, x10_c, x11, x12_c, x13, x14, x15, x16, x17_c, x18, x19_c, x20, x21, x22, x24, x25_c, x26_c, x27, x28, x30, x31, x32, x34_c, x36_c, x37_c, x38_c, x39_c, x40, x41_c, x42_c, x44, x45, x46, x47_c, x48, x50_c, x51_c, x52_c, x53, x54_c, x56_c, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75, x76_c, x79_c, x80_c, x81_c, x82, x83, x84, x85_c, x86, x87_c, x88_c, x89_c, x91, x92_c, x94_c, x95_c, x96, x97_c, x99);
and (w19, x5_c, x6, x7, x8, x9_c, x12_c, x14, x16_c, x17_c, x18, x19, x22_c, x23_c, x26, x30, x31_c, x33, x34, x36, x40, x47_c, x48, x53, x54_c, x57_c, x58, x61_c, x62, x65_c, x66, x68_c, x69_c, x70, x71, x72, x73_c, x75_c, x81_c, x86_c, x88, x89_c, x91, x92_c, x93_c, x98_c);
and (w20, x15, x20, x21_c, x29, x41, x49_c, x58, x63_c, x64, x70, x99);
and (w21, x5_c, x8_c, x9, x11, x12_c, x13, x14_c, x15_c, x16_c, x19_c, x21_c, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37, x38, x40, x45, x46_c, x47, x49, x50, x51_c, x55_c, x56, x57_c, x58, x59_c, x60, x62, x64, x65_c, x66, x68_c, x69_c, x70_c, x71, x72_c, x74_c, x76_c, x77, x78_c, x81, x85, x87_c, x88, x90, x91, x93, x94_c, x95, x97_c, x98_c, x99_c);
assign w22 = x94;
and (w23, x3_c, x8, x13_c, x15, x17_c, x27, x28_c, x29, x31_c, x38_c, x40, x42, x43_c, x44_c, x46_c, x49, x52_c, x53, x56_c, x57_c, x58_c, x60, x63_c, x69, x75_c, x76_c, x77_c, x79, x84, x85_c, x92_c, x98);
and (w24, x1, x3_c, x4_c, x6, x7, x8, x10_c, x12, x13, x14_c, x16, x18_c, x20_c, x22, x23, x24_c, x26_c, x27, x29, x33, x34_c, x35, x36_c, x39, x41, x42, x43, x46_c, x48, x53, x54, x56, x57, x58, x61, x62_c, x63, x64, x68_c, x71_c, x73, x76_c, x77_c, x78_c, x80, x86_c, x89, x93_c, x99);
and (w25, x0, x1, x2_c, x3_c, x4_c, x5, x6_c, x8_c, x10_c, x11, x12, x13, x14, x15_c, x16, x18_c, x19_c, x20, x21_c, x22_c, x26_c, x27_c, x28_c, x29_c, x31, x32, x33, x34_c, x36, x37_c, x38_c, x39_c, x40, x41, x42, x43, x44, x46_c, x47, x49, x50_c, x52_c, x53, x54, x55_c, x56_c, x57_c, x58, x59_c, x61_c, x62_c, x63, x64_c, x66_c, x67_c, x68_c, x73, x75_c, x76, x77_c, x78_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x86_c, x87_c, x88_c, x89, x90, x91_c, x92, x96_c, x97, x98_c);
and (w26, x1_c, x2, x3_c, x4, x11_c, x12, x14, x15, x16, x18_c, x20, x21_c, x22_c, x24, x26_c, x27_c, x29, x30_c, x32_c, x33_c, x34_c, x35, x36, x37_c, x40, x43, x44, x47, x50_c, x52_c, x53_c, x54_c, x55_c, x56_c, x58, x59_c, x60, x63, x69, x70, x73_c, x76, x77_c, x82_c, x83_c, x84, x88, x89_c, x90, x92, x95, x97_c, x98_c);
and (w27, x0, x1, x2_c, x3, x4, x5, x6_c, x7, x9, x10_c, x11_c, x12_c, x13_c, x14, x15, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23, x24, x25, x26_c, x27, x28_c, x29_c, x30, x31, x32, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40, x41, x42_c, x43_c, x44, x45, x46, x47_c, x48, x49, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67, x68, x69_c, x70_c, x71, x72, x73, x74, x75, x76_c, x77, x79_c, x80_c, x81_c, x83_c, x84_c, x85, x87, x88, x89_c, x90_c, x91_c, x92_c, x93, x94, x95_c, x96_c, x97, x98_c, x99);
and (w28, x2_c, x4_c, x5, x6_c, x9, x10_c, x12_c, x16, x18, x19, x20_c, x21_c, x22, x24, x25_c, x26, x27_c, x28, x31, x32_c, x33, x34, x36, x37, x38_c, x39, x40_c, x41, x44, x45, x46_c, x47_c, x48, x49, x50, x51, x52, x53_c, x54, x56, x57_c, x58_c, x60, x61_c, x62, x64_c, x65_c, x66, x67_c, x70, x71, x72_c, x74, x76, x80, x81_c, x83, x85, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93, x98, x99);
and (w29, x18_c, x24, x25_c, x26, x28_c, x30, x31_c, x34_c, x36, x42_c, x48_c, x51_c, x53, x56_c, x59_c, x79_c, x80, x81_c, x83, x92_c, x94, x95, x99_c);
and (w30, x0_c, x2_c, x3, x4_c, x6_c, x15, x16_c, x17, x21, x23, x26, x28, x30_c, x31, x32, x35_c, x36, x37_c, x38, x39_c, x41, x43_c, x46_c, x47_c, x49, x51_c, x56_c, x59, x63_c, x64, x65, x68, x70, x75_c, x76_c, x81_c, x82, x84, x87_c, x88, x89, x90_c, x92, x99_c);
and (w31, x0_c, x4_c, x7, x8, x11, x12, x14, x18_c, x21, x25, x30_c, x31_c, x38, x41, x43_c, x44_c, x45, x50, x52, x55_c, x58, x60_c, x68_c, x69_c, x70_c, x71_c, x74, x76_c, x77, x85, x89_c, x90, x93_c, x99_c);
and (w32, x3_c, x4, x5, x6, x7_c, x9, x12_c, x13, x14, x15, x18, x24_c, x27_c, x31, x32, x34, x36_c, x38, x40_c, x44, x48_c, x49, x53, x56_c, x57, x58, x59, x60, x61, x62, x65, x66_c, x67, x70, x71_c, x73_c, x75_c, x76_c, x78, x81, x83, x85, x87_c, x88_c, x94, x95, x96_c);
and (w33, x0, x1, x5_c, x11_c, x14, x26, x31_c, x32_c, x34_c, x35, x36_c, x37_c, x38, x45_c, x51, x52_c, x53_c, x54_c, x62_c, x63, x72_c, x76, x77, x81, x82, x83_c, x85, x86_c, x88_c, x92, x94, x98_c);
and (w34, x3_c, x6_c, x8_c, x11_c, x12_c, x16_c, x18, x21, x23, x25_c, x32, x33, x34_c, x36, x43_c, x46, x52, x53, x58, x59_c, x60, x62_c, x64, x66_c, x71_c, x72_c, x79, x80, x81_c, x88_c, x90_c, x92, x98_c);
and (w35, x8_c, x14_c, x23, x26, x38, x51_c, x62_c, x70, x77_c, x92_c, x99_c);
and (w36, x0, x4, x5_c, x6, x7, x9, x11_c, x12_c, x13_c, x15_c, x16, x18_c, x19, x20, x23_c, x25_c, x26_c, x27_c, x28, x30, x31, x33_c, x35, x39_c, x40_c, x42, x44_c, x48, x49, x50, x51, x53, x54, x57_c, x58, x60, x61_c, x65_c, x66_c, x68, x70, x73, x74, x76_c, x79_c, x80, x81_c, x82, x83_c, x85_c, x86, x87, x88_c, x90, x91_c, x92, x95, x97);
and (w37, x2_c, x4, x5, x6_c, x11_c, x13, x16, x21, x23, x31, x32_c, x33_c, x34, x36, x38_c, x40, x43_c, x46_c, x47, x48_c, x50_c, x56_c, x61, x62_c, x65_c, x67, x68_c, x73_c, x74_c, x77_c, x78, x80_c, x82, x83, x85, x88_c, x89_c, x90_c, x92, x93, x95, x96_c, x97_c);
and (w38, x1_c, x4_c, x5, x16, x22_c, x28, x29_c, x33, x38, x41, x42_c, x49_c, x56, x67, x75_c, x81_c, x84_c, x88_c, x91, x94_c, x98_c);
and (w39, x0_c, x1_c, x2, x3_c, x6, x7, x8_c, x9_c, x12_c, x13, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x23_c, x24, x25, x26, x27, x28, x30, x31_c, x32, x34, x35_c, x36_c, x37, x38_c, x39, x41_c, x42_c, x43_c, x44, x45_c, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x55_c, x56, x57_c, x58_c, x59, x61, x62_c, x63, x64_c, x65_c, x66_c, x67, x68, x69_c, x70, x71_c, x72, x73, x74, x75, x76, x77, x78, x80_c, x83_c, x84, x85_c, x86, x87_c, x88, x89_c, x90_c, x93_c, x94, x96, x97, x98_c, x99_c);
and (w40, x0, x4, x5, x6, x8, x9, x11, x12, x13, x15_c, x16, x17, x18_c, x19, x23_c, x24_c, x26_c, x27, x28_c, x29_c, x31, x35, x37, x38_c, x39_c, x40, x41, x42_c, x43_c, x44_c, x49_c, x52, x53_c, x54, x56, x57_c, x62, x63_c, x65_c, x66_c, x69, x70, x72_c, x74, x76, x78, x79, x80, x83_c, x85, x86_c, x88_c, x91_c, x92, x95_c, x96_c, x97_c, x98);
and (w41, x11, x21, x27, x33_c, x53_c, x60, x72_c, x84_c, x85_c, x87);
and (w42, x0_c, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21, x22_c, x24, x25_c, x27_c, x28_c, x29, x30, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46, x47, x48, x49, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x62_c, x65_c, x66, x67, x68_c, x69, x71_c, x72, x74_c, x76, x79, x80_c, x81_c, x82_c, x84, x85, x86, x87_c, x88_c, x89, x91, x93_c, x94_c, x95_c, x96, x97, x98, x99_c);
and (w43, x0_c, x1, x2_c, x4, x5, x9_c, x10_c, x12_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19, x20_c, x21_c, x22_c, x24, x25_c, x26_c, x28, x29, x30_c, x32, x33_c, x34, x35, x36_c, x37_c, x38, x39, x40, x42, x43, x44, x45_c, x46, x47, x48_c, x50_c, x51_c, x52, x53_c, x55_c, x56, x57, x59, x60_c, x62, x63_c, x64, x66, x67_c, x68, x69_c, x71, x72_c, x73, x74_c, x75_c, x76_c, x78_c, x81_c, x83_c, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93, x95_c, x96, x97_c, x98_c, x99);
and (w44, x0_c, x3, x5_c, x10_c, x14_c, x19, x25, x26_c, x29, x30_c, x33_c, x37, x39_c, x42_c, x43, x44_c, x49_c, x51, x61, x64_c, x67_c, x68, x69_c, x72, x78_c, x92_c, x97_c, x99);
and (w45, x7_c, x8, x15_c, x18_c, x19, x20, x23_c, x25_c, x36, x44_c, x51_c, x57, x59_c, x62, x64_c, x70, x74, x79, x80, x81_c, x90_c, x91_c, x97_c, x99_c);
and (w46, x1_c, x2, x3_c, x4, x5, x6_c, x7_c, x8, x9_c, x11, x12_c, x13, x14_c, x15, x16_c, x17_c, x18_c, x19_c, x20, x21, x23, x24_c, x25_c, x26, x27, x28, x29, x30_c, x31_c, x32, x33_c, x34, x35_c, x36_c, x38, x39_c, x40_c, x41_c, x42, x43, x44_c, x45, x46_c, x47, x48, x49, x50, x51, x52_c, x53, x54, x55_c, x56_c, x57_c, x58_c, x60, x61, x62, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x73, x74, x75, x76_c, x77_c, x78, x79, x80_c, x81_c, x82, x83, x84, x85_c, x86, x87, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97, x98_c, x99_c);
and (w47, x4, x6, x7_c, x8, x10_c, x16_c, x29, x35, x36, x38_c, x45, x51, x53, x54_c, x56, x57, x66, x69, x72_c, x73_c, x74, x76, x78, x79, x82_c, x83, x84_c, x85, x86_c, x88, x92_c);
and (w48, x1, x2, x5_c, x7, x12_c, x16_c, x19, x26, x30, x31, x32_c, x36, x38_c, x40_c, x42_c, x43_c, x48_c, x49_c, x56_c, x60_c, x62_c, x65_c, x70_c, x73_c, x75_c, x79, x81_c, x84_c, x85, x87_c, x88, x91_c, x93_c, x94, x98_c);
and (w49, x3, x5, x7, x12_c, x21_c, x25, x28, x35, x39, x41, x47, x48, x56, x57_c, x59, x65_c, x68_c, x71, x76_c, x79_c, x81, x88_c, x89, x90_c, x95_c, x97_c, x98, x99_c);
and (w50, x16, x38, x55, x63, x77, x82_c, x93);
and (w51, x0, x1, x2, x3_c, x5_c, x8_c, x9, x10_c, x14, x16, x17, x18, x21_c, x22, x24, x25_c, x26, x30_c, x31, x32, x33, x34_c, x36, x38_c, x39_c, x40, x41_c, x42_c, x45, x46, x47, x48_c, x49, x50, x51, x53, x54, x55, x57, x60, x61, x62, x64_c, x66_c, x69, x70_c, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80, x81, x82_c, x83, x90, x91, x92, x93_c, x94, x96_c, x97, x99);
and (w52, x2, x3, x5_c, x6_c, x10, x11, x12_c, x13, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x23_c, x24_c, x26, x28, x31_c, x32, x33_c, x34, x38, x39_c, x41_c, x43, x44_c, x45_c, x46_c, x47, x51_c, x52, x54, x62_c, x65, x66_c, x67_c, x68, x71, x73_c, x75_c, x77, x79, x80_c, x81, x82, x84, x85_c, x86_c, x87_c, x89_c, x90, x91, x92, x94, x96, x97_c, x98_c);
and (w53, x0, x1_c, x2_c, x4_c, x5, x16, x17, x18, x19, x20_c, x21_c, x22_c, x24_c, x25, x27_c, x28_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x36_c, x38, x40_c, x43, x44, x45, x46, x47, x51_c, x52_c, x53_c, x54, x56_c, x58_c, x61, x62, x64_c, x65, x66, x68_c, x71_c, x72, x73, x74_c, x76_c, x77, x81, x87, x89, x91, x94_c, x95_c, x96, x99);
and (w54, x1, x2_c, x3_c, x5_c, x6_c, x7, x10_c, x12_c, x13_c, x14_c, x15, x16_c, x17, x21_c, x22_c, x25, x26, x27_c, x32_c, x34_c, x36, x38, x40_c, x41_c, x42, x43, x45, x46_c, x48_c, x49, x50, x51_c, x52, x53, x55, x57, x58, x61_c, x62, x64_c, x65_c, x66, x67_c, x68_c, x69_c, x70, x76_c, x77, x78, x79_c, x80, x81, x82_c, x84, x85_c, x87, x88_c, x89_c, x93, x94, x96_c, x99_c);
and (w55, x0_c, x1_c, x2, x6, x7_c, x8, x10, x11, x12_c, x13, x14_c, x15, x17_c, x18, x19_c, x20_c, x21, x22_c, x24, x25, x26, x28, x29, x30, x31_c, x32_c, x33_c, x34_c, x36_c, x37_c, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49, x51_c, x52_c, x53_c, x54, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x69, x71_c, x72_c, x73, x75, x76_c, x77, x79_c, x80_c, x81, x83_c, x84_c, x85, x86_c, x87_c, x88_c, x89, x90, x91_c, x92, x93, x94, x95, x96_c, x97, x98_c, x99_c);
and (w56, x0, x2, x4_c, x6, x7_c, x9_c, x13_c, x15, x16, x19, x20, x24, x27, x29_c, x31_c, x33_c, x35, x37_c, x38_c, x39, x45_c, x50_c, x51, x52_c, x55_c, x56, x59_c, x61_c, x73_c, x76_c, x82, x89, x92_c, x95, x96_c);
and (w57, x0_c, x1_c, x2, x3_c, x4, x5_c, x6_c, x7_c, x8, x9, x10, x11_c, x12_c, x13, x14_c, x15, x16_c, x17_c, x18, x19_c, x20, x21_c, x22_c, x23_c, x24_c, x25, x27_c, x28, x29, x30_c, x31, x32_c, x33, x34, x36_c, x37, x38, x39_c, x40, x41_c, x42, x43, x44, x45, x46_c, x47_c, x48_c, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56, x57_c, x58_c, x59_c, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x67, x68_c, x69, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80, x81_c, x82_c, x83, x84, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91, x92_c, x93, x94, x95, x96, x97, x98_c, x99_c);
and (w58, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x11_c, x12, x13, x15_c, x16_c, x17_c, x18, x19, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x27_c, x29, x30, x31, x32, x34_c, x36, x37_c, x38_c, x41, x42_c, x43_c, x44, x46, x49_c, x51, x53, x55, x56_c, x57, x58, x59_c, x60, x61_c, x64, x65, x66_c, x67_c, x70, x71, x72_c, x73_c, x74, x75, x76_c, x77, x78_c, x79, x80, x82_c, x83_c, x84_c, x85_c, x86, x87, x88, x89, x90, x92, x96_c, x97);
and (w59, x0_c, x6_c, x9, x11_c, x19, x23_c, x26, x32, x35_c, x45_c, x48, x55, x57, x58_c, x61, x67_c, x69_c, x71, x75, x77, x80, x84_c, x85_c, x87_c, x91_c, x96_c, x97_c, x98);
and (w60, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7, x8, x9_c, x10, x11_c, x12_c, x13, x14, x16_c, x17_c, x18, x19, x20_c, x21, x22, x23, x24_c, x26, x27_c, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x41_c, x42, x43, x44, x45, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55_c, x56, x57_c, x59_c, x60_c, x61, x62, x63_c, x64_c, x65, x66, x67_c, x68, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x76_c, x77_c, x78, x79_c, x80, x81_c, x82, x83, x84_c, x86, x87, x88, x89, x90, x91, x92_c, x93_c, x94, x95_c, x96, x97, x98_c);
and (w61, x0, x1, x2_c, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12, x13_c, x14, x15, x16_c, x17_c, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x28, x29, x30_c, x31_c, x32, x33_c, x34_c, x35_c, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x45, x46, x47_c, x48, x49_c, x50, x51_c, x52_c, x53, x54, x55_c, x56, x57, x58_c, x59_c, x60_c, x61, x62, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73, x74, x75_c, x76_c, x77, x78_c, x79_c, x81_c, x82_c, x83, x85_c, x86, x87, x88, x89_c, x90, x91, x92_c, x93, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w62, x3, x7_c, x8_c, x13_c, x17_c, x19, x21_c, x26, x29, x38_c, x39, x42, x45, x47, x57, x62, x75_c, x80_c, x81, x86, x90, x93, x94, x96_c, x97, x99_c);
and (w63, x0, x1_c, x4, x5, x6_c, x7, x8, x9, x11, x12_c, x13_c, x15_c, x16, x18_c, x20, x21, x22, x23, x24, x25, x26_c, x29_c, x30, x31_c, x32, x33_c, x35_c, x36_c, x37_c, x38, x39, x40, x41_c, x44_c, x45, x46, x47, x49, x50_c, x51, x52_c, x53_c, x54_c, x55_c, x56, x57_c, x58, x59, x60, x61, x63, x64, x65, x66, x68_c, x69, x70, x71, x74_c, x76_c, x78, x80_c, x81_c, x82, x83_c, x85, x90_c, x92_c, x93, x94_c, x96_c, x98);
and (w64, x2, x9, x11, x15, x16, x17_c, x18_c, x19_c, x23, x24_c, x25, x27_c, x28_c, x29, x30, x35, x36_c, x39, x40_c, x41_c, x44_c, x47, x48_c, x51, x55_c, x58, x68, x70_c, x73_c, x74_c, x75, x76, x77_c, x78, x81, x82_c, x83_c, x86_c, x88, x89_c, x95, x96_c, x97_c);
and (w65, x16_c, x26_c, x34_c, x45, x73_c, x75_c, x78_c, x79, x81, x83_c, x88, x91_c);
and (w66, x0_c, x2, x3_c, x4, x5, x6, x7_c, x9_c, x10_c, x13, x14, x15, x17_c, x18, x19, x21_c, x23, x24, x25_c, x26_c, x27, x29_c, x30, x32, x33_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41, x42, x43, x44_c, x45, x46, x47, x48_c, x50, x51, x52, x53_c, x54_c, x55, x58, x59_c, x60_c, x61_c, x62, x63, x64, x65_c, x66_c, x67_c, x68_c, x70_c, x71_c, x73_c, x74_c, x75_c, x77_c, x78, x79, x80_c, x81_c, x82, x83_c, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91, x94, x95, x97_c, x98, x99);
assign w67 = x52_c;
and (w68, x0, x1, x2_c, x3_c, x4, x5, x6, x7, x8, x9, x10_c, x11, x12_c, x13_c, x14_c, x15, x16_c, x17, x18_c, x19_c, x20_c, x21, x22, x23, x24_c, x25, x26, x27_c, x28, x29, x30_c, x31_c, x32_c, x33, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x44_c, x45, x46_c, x47, x48_c, x49_c, x50_c, x51_c, x52, x53, x54_c, x56, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x66, x67_c, x68, x69_c, x70_c, x71, x72, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x84, x85_c, x86, x87_c, x88_c, x89, x90, x91_c, x92, x93_c, x94_c, x95_c, x96, x97_c, x98_c, x99_c);
and (w69, x3_c, x8, x12, x19_c, x23_c, x33, x36_c, x42_c, x46_c, x55_c, x56, x59, x61, x64_c, x67, x71, x74, x77, x78_c, x84_c, x88, x93_c);
and (w70, x0, x1, x2, x3_c, x5_c, x6_c, x7_c, x8_c, x9, x10, x11_c, x12_c, x14, x15_c, x16_c, x17_c, x18, x19, x20, x21, x22, x23, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31_c, x32_c, x33, x34_c, x35, x36_c, x37_c, x38, x39, x40, x41, x42, x43, x44_c, x45, x46_c, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54, x55_c, x56_c, x57_c, x58_c, x59_c, x60, x61, x62_c, x63, x64_c, x65, x66, x67, x68_c, x69_c, x70, x72_c, x73_c, x74, x75_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99_c);
and (w71, x3_c, x9, x10_c, x13, x16, x17, x19, x20, x21, x25_c, x28, x30, x34_c, x35, x39, x41_c, x44_c, x46_c, x48, x50, x54, x55, x60_c, x61_c, x62_c, x63, x65, x67_c, x68_c, x70, x71_c, x73, x75, x78, x79_c, x81_c, x82, x83_c, x87_c, x89_c, x93_c, x97_c);
and (w72, x3, x9_c, x11_c, x19, x24_c, x27_c, x35_c, x39, x55, x56_c, x72, x89_c);
and (w73, x0, x1, x2, x3_c, x4_c, x5_c, x6, x7_c, x8, x9, x10, x11, x12_c, x13, x14, x15, x16, x17, x18, x19_c, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x27, x28, x29, x30_c, x31, x32_c, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45, x46_c, x47, x48_c, x49_c, x50_c, x51, x52, x53_c, x54_c, x55_c, x56, x57, x58, x59_c, x60_c, x61, x62, x63_c, x64_c, x65, x66, x67, x68_c, x69, x70, x71_c, x72, x73_c, x74, x75, x76, x77, x78, x79_c, x80_c, x81, x82, x83, x84, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w74, x2, x4_c, x5, x6, x7_c, x9_c, x13, x16_c, x17, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x25, x27, x28, x31_c, x33_c, x34, x36, x39, x41, x42, x43, x45_c, x47_c, x48_c, x49_c, x51, x52, x53_c, x54_c, x56_c, x57_c, x58_c, x59, x62, x63_c, x65, x67_c, x68_c, x71_c, x72_c, x73, x74, x75, x78, x80, x81, x82_c, x84_c, x86, x87, x88_c, x89, x90_c, x92_c, x94, x96_c, x97);
and (w75, x0_c, x1, x2, x5_c, x6, x7_c, x10, x13_c, x14, x16, x17_c, x22, x24_c, x26, x29, x30_c, x32, x35, x37, x38_c, x39_c, x40_c, x43_c, x44_c, x45_c, x47, x48_c, x50, x54_c, x56_c, x58_c, x59, x60_c, x61_c, x62, x65, x67, x68, x71, x73_c, x76_c, x80_c, x81, x83_c, x84, x85_c, x88, x89_c, x90_c, x92_c, x96);
and (w76, x0, x2_c, x4_c, x6, x7, x9_c, x10, x11, x13_c, x15, x17, x18, x19, x20, x22, x23, x25, x26_c, x28, x29_c, x31_c, x33_c, x35_c, x36_c, x37_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x46, x49_c, x51, x52, x55_c, x58_c, x60, x65_c, x66, x67_c, x69, x70_c, x71, x73, x74, x75, x78, x80_c, x81, x82, x84_c, x86_c, x87, x89, x91, x94, x96_c);
and (w77, x0, x3, x5, x6, x9, x10, x11_c, x14, x15_c, x18_c, x20, x21, x25_c, x26_c, x27_c, x28_c, x29, x31, x37_c, x38_c, x39_c, x42_c, x43, x44_c, x50, x51_c, x52, x53_c, x57, x58, x62_c, x63, x64, x67_c, x69, x71_c, x73_c, x74, x75_c, x81_c, x82, x83_c, x86_c, x87, x88_c, x89, x90, x92_c, x96_c, x97_c);
and (w78, x0, x2, x3_c, x4, x5_c, x7, x8, x9, x13_c, x18_c, x20, x27_c, x29, x30_c, x31, x34, x36_c, x40_c, x42, x43, x47_c, x50, x51, x53, x54, x55, x57_c, x59, x62, x65_c, x66, x71, x75, x77_c, x79_c, x80_c, x81_c, x82_c, x83_c, x84, x87_c, x89);
and (w79, x0_c, x1, x2_c, x7_c, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14_c, x15, x16, x18, x19, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26, x27, x29, x30, x31_c, x34, x35, x36, x37, x38_c, x40_c, x41, x42, x44_c, x45_c, x46_c, x48, x49, x50_c, x51_c, x53, x54, x55, x56_c, x57, x58_c, x59, x60, x62_c, x64_c, x65, x66, x67_c, x68_c, x70, x71, x72_c, x73_c, x74, x75_c, x76_c, x77, x80_c, x81, x83_c, x84, x85, x86, x87, x90, x91, x92_c, x93_c, x94, x95_c, x98, x99_c);
and (w80, x0_c, x1, x3_c, x5_c, x6, x7, x8, x9, x10, x11_c, x12_c, x14, x15_c, x16, x17_c, x18, x20_c, x21, x22, x23_c, x25, x26_c, x27, x28_c, x31_c, x32, x33, x35_c, x36_c, x37, x38_c, x39, x42, x46_c, x47_c, x49_c, x51_c, x52_c, x53_c, x54, x55, x56_c, x57, x59_c, x60_c, x62, x63_c, x64, x66, x69_c, x70_c, x71, x72_c, x75, x77_c, x80_c, x81_c, x82_c, x84, x85_c, x86_c, x87_c, x89, x90, x91_c, x93, x94, x99_c);
and (w81, x2, x5, x6_c, x8_c, x9_c, x13_c, x14_c, x15_c, x16, x17, x18_c, x22, x23_c, x24_c, x28_c, x29, x30_c, x31_c, x34, x35, x36_c, x37, x38_c, x39, x40_c, x41_c, x42, x44_c, x45_c, x46_c, x47_c, x49, x51_c, x54, x55_c, x56_c, x57, x58, x59_c, x60_c, x62_c, x64, x65_c, x66_c, x69, x72_c, x74, x75_c, x79, x80_c, x82, x83, x85, x87, x88, x89, x90_c, x92, x93_c, x95, x97_c, x98, x99);
and (w82, x0, x1, x2_c, x5_c, x7, x8_c, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18_c, x19_c, x20, x21_c, x22, x23, x24, x26_c, x27_c, x29_c, x30_c, x31, x32_c, x34_c, x35_c, x36, x37_c, x38_c, x40, x42_c, x43_c, x44_c, x45, x46, x47, x48_c, x49, x51_c, x52_c, x53, x54, x55_c, x56_c, x57, x58_c, x59_c, x60_c, x61_c, x62_c, x63_c, x64, x65, x66_c, x67, x68_c, x69, x70_c, x71_c, x72, x73, x74, x75, x76, x77, x78_c, x79_c, x82_c, x83, x84, x85, x86_c, x87, x88, x89, x90, x91, x94_c, x95_c, x96, x97_c);
and (w83, x4_c, x14_c);
and (w84, x0_c, x1, x2, x4, x14, x16, x17_c, x20_c, x22_c, x23_c, x25, x31_c, x33_c, x38_c, x44, x45_c, x47, x53, x54_c, x55, x56_c, x57_c, x61_c, x63_c, x70_c, x74, x78_c, x83_c, x84, x85_c, x86, x90_c, x92_c, x94_c, x95, x96, x97, x99);
and (w85, x2_c, x3_c, x4_c, x6, x7, x8, x10_c, x12, x13, x16, x17_c, x18, x20_c, x21_c, x25_c, x26, x28_c, x36_c, x38_c, x39, x40, x41_c, x42_c, x43, x45, x46, x47_c, x61_c, x66, x70_c, x74_c, x76, x80, x81_c, x82_c, x83_c, x84_c, x87, x88_c, x90, x94_c, x97_c, x98);
and (w86, x2_c, x3, x4, x6_c, x11_c, x13_c, x14, x15_c, x18_c, x19_c, x20_c, x22_c, x23, x25, x27, x29_c, x30, x32_c, x33_c, x34_c, x39_c, x40, x43, x44_c, x47_c, x49, x50_c, x52, x53, x56, x60, x62_c, x66, x67, x68_c, x72_c, x73_c, x74_c, x75, x77_c, x78, x80, x81, x82, x84_c, x85_c, x86, x87, x90, x93, x95, x96_c, x97_c);
assign w87 = x19;
and (w88, x4_c, x9_c, x14, x16_c, x25_c, x34_c, x55_c, x61, x75_c, x76, x83_c, x86_c, x88, x89_c);
and (w89, x9, x12, x13_c, x14_c, x23_c, x31_c, x32_c, x43_c, x45_c, x48, x51_c, x52_c, x54, x55, x68, x87_c, x94, x95, x96_c);
and (w90, x0_c, x2, x3, x4_c, x5, x8_c, x10, x11, x12, x13, x14_c, x15_c, x17_c, x18, x19_c, x20, x21, x22, x23, x24_c, x25_c, x27_c, x29, x30_c, x31, x33, x34, x35, x36, x37, x38, x40_c, x41_c, x42, x43, x44_c, x45, x46_c, x47_c, x49_c, x50, x52_c, x53, x54_c, x55, x56, x57_c, x58_c, x61_c, x62, x63, x65_c, x66, x67, x68, x69, x70, x72, x73, x74_c, x75, x76_c, x78_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x87_c, x88_c, x90, x91, x92_c, x93, x94, x95_c, x97);
and (w91, x0, x1, x2_c, x4, x5_c, x6, x7_c, x8, x9, x10, x11, x13, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x30, x31_c, x32, x33_c, x34, x35, x36_c, x37, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46, x47_c, x48, x49_c, x50_c, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62_c, x63_c, x64, x65_c, x66, x67_c, x68_c, x69_c, x70, x71, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x79, x80, x81_c, x82, x83_c, x84, x86, x87, x88, x89, x90_c, x91, x92, x93, x94_c, x95, x96, x97, x98_c, x99);
and (w92, x0, x2_c, x3_c, x4, x6_c, x7, x8, x11, x12, x13, x14, x17, x19_c, x20_c, x21_c, x22_c, x23_c, x24, x25, x27, x28_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x37_c, x38_c, x41_c, x42_c, x43, x44, x46, x47_c, x50, x54, x55_c, x56_c, x57_c, x58_c, x59_c, x61, x62_c, x63_c, x64_c, x66, x67_c, x68, x69_c, x70_c, x71_c, x72, x73_c, x74_c, x75_c, x77_c, x78, x79_c, x80, x82, x83, x84_c, x85_c, x86, x87_c, x88, x90_c, x91_c, x95, x96, x98_c, x99);
and (w93, x2, x3_c, x4, x6, x9, x10_c, x11_c, x12, x18, x19_c, x21_c, x22, x23, x25, x26, x30_c, x34_c, x35, x39_c, x40_c, x42_c, x43_c, x45, x47_c, x54_c, x58_c, x59, x63_c, x66_c, x67_c, x69_c, x70, x72, x78_c, x81, x83, x84_c, x85_c, x86_c, x94, x95_c, x98_c);
and (w94, x0, x1_c, x2, x3, x5_c, x6_c, x7, x8_c, x9_c, x10_c, x11, x12, x14, x16_c, x17, x18, x19, x20_c, x21_c, x22_c, x23_c, x25_c, x26_c, x27, x28, x29_c, x30, x31, x32_c, x33, x34, x35_c, x36, x37, x38, x39_c, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x52_c, x53_c, x54, x55_c, x58_c, x59_c, x60, x61, x62, x63, x65, x66_c, x67_c, x69, x70, x71, x72_c, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84, x85, x86, x87, x88, x89_c, x90_c, x91_c, x92, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w95, x0, x1_c, x2, x3, x4_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12_c, x16, x18, x19, x20_c, x22_c, x25, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36, x37, x38_c, x39, x40, x42_c, x44, x45_c, x46, x47, x48, x49, x50, x52_c, x54, x55_c, x58_c, x59_c, x60_c, x61_c, x62_c, x64, x65_c, x66, x67, x68_c, x71_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81_c, x83_c, x84_c, x86, x88, x89_c, x91, x93, x95, x96, x97, x98_c, x99);
and (w96, x21, x22, x23_c, x27_c, x68, x81_c, x83, x94_c, x98);
and (w97, x0_c, x1, x2, x3, x4, x5, x6, x7, x8_c, x9, x10_c, x11, x12, x14, x15, x16, x17_c, x18, x19, x21_c, x22, x23, x24_c, x25_c, x26, x27_c, x28_c, x31, x32_c, x33, x34, x35, x36, x37_c, x38, x40_c, x41_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x52, x53_c, x56_c, x57, x58, x59_c, x60, x61_c, x62_c, x63, x64, x66_c, x67_c, x68_c, x70, x71_c, x72, x73, x75, x78, x79_c, x81, x82_c, x83, x84, x85_c, x86, x88_c, x89_c, x90_c, x91_c, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w98, x3, x5_c, x18, x21_c, x33_c, x39_c, x76, x77_c, x94);
and (w99, x4_c, x27, x28, x34_c, x36, x41, x53, x54_c, x57_c, x66, x68_c);
and (w100, x0_c, x1_c, x3, x4_c, x6, x7_c, x8, x10_c, x12, x13, x14, x18, x19, x20, x21_c, x24_c, x25, x27, x28, x29, x30, x31_c, x32_c, x34, x37, x38_c, x39, x41_c, x44, x49_c, x54_c, x56_c, x59_c, x60, x62, x63, x64_c, x65_c, x66, x67_c, x68_c, x70, x71_c, x73, x74_c, x76_c, x77, x78_c, x82, x85, x90, x91, x93, x94, x96, x97);
and (w101, x0, x1_c, x2_c, x3, x4_c, x5_c, x6_c, x7_c, x9_c, x10_c, x11, x12_c, x13, x14_c, x15_c, x17_c, x18_c, x19, x20_c, x21, x22, x23, x24_c, x25, x26, x27_c, x28_c, x29, x30_c, x31, x32_c, x33, x34, x35_c, x37_c, x38_c, x39, x40_c, x41_c, x42, x43_c, x44_c, x46, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54, x55_c, x56_c, x57, x58_c, x59, x60_c, x61_c, x62_c, x63, x64, x65, x66, x67_c, x68, x70, x71, x72, x73_c, x74, x75_c, x76, x77_c, x78, x79_c, x80, x81, x82, x83_c, x84, x85, x86_c, x87, x88_c, x89, x90_c, x91_c, x92_c, x93, x95_c, x96_c, x97_c, x98, x99);
and (w102, x0_c, x2, x3_c, x8_c, x12, x22, x24_c, x28_c, x29_c, x33, x35, x39, x40_c, x46_c, x48, x53_c, x55_c, x60_c, x66, x72, x75_c, x78, x82, x83, x86, x87, x95, x96_c, x97_c);
and (w103, x1, x4_c, x10_c, x11_c, x13_c, x14, x15_c, x19_c, x22, x24, x25_c, x28_c, x31, x35_c, x36_c, x39_c, x41_c, x45, x50, x54, x62, x63, x64, x66_c, x72_c, x76_c, x77, x82, x87, x90, x96_c, x99_c);
and (w104, x0_c, x1, x2_c, x5, x6_c, x7_c, x9_c, x10, x11, x12_c, x13, x14, x15, x16_c, x17, x19_c, x20, x21_c, x22_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x36_c, x37, x38, x39_c, x40, x41_c, x42, x43_c, x44_c, x45_c, x46, x47, x48_c, x49_c, x50_c, x52_c, x53_c, x54_c, x55, x56, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x76, x77, x78_c, x79_c, x80_c, x81_c, x82, x83, x84_c, x85_c, x86, x87_c, x89, x90, x91, x92_c, x93, x94, x95_c, x96_c, x98_c, x99);
and (w105, x7_c, x9_c, x13, x14, x21, x45_c, x50_c, x59, x61_c, x63_c, x65_c, x72, x77_c, x78, x79, x83, x84, x89_c);
and (w106, x0, x1, x2, x3_c, x4, x5, x6, x7, x8, x9, x10_c, x11, x12_c, x13, x14_c, x15_c, x16, x17, x18_c, x19_c, x20, x21_c, x22_c, x23, x25_c, x26_c, x27_c, x28_c, x29, x30_c, x31, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x40_c, x41_c, x43, x44, x45_c, x48_c, x50_c, x51_c, x52, x53, x54, x55_c, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x67_c, x68, x69_c, x70_c, x71, x72_c, x73, x74_c, x76_c, x77_c, x78_c, x79, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x89, x90_c, x91, x93_c, x94_c, x95, x96_c, x97, x98_c, x99);
and (w107, x3_c, x7, x8_c, x19_c, x30_c, x34, x38_c, x55_c, x61_c, x68, x69, x72, x77, x78, x85_c, x87, x89_c, x94, x95_c, x98);
and (w108, x0_c, x1_c, x2_c, x3, x4_c, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13, x14_c, x15_c, x16, x17, x18_c, x19_c, x20, x21, x22_c, x23, x24_c, x25_c, x26, x27_c, x28_c, x29, x30_c, x31_c, x33_c, x34_c, x35_c, x36_c, x37_c, x38, x39_c, x41_c, x42, x43_c, x44, x46_c, x47, x48_c, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56, x57_c, x58_c, x59, x60_c, x61_c, x62, x63_c, x64_c, x65, x66_c, x67, x68, x69, x70_c, x72_c, x73, x74, x75, x76, x77, x78_c, x79_c, x80_c, x82_c, x83, x84_c, x85_c, x86_c, x87, x88, x90_c, x91, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w109, x0_c, x2_c, x3_c, x6, x7_c, x10, x11, x14_c, x15_c, x16, x17, x21_c, x23_c, x25, x27, x28_c, x29, x30, x31_c, x32, x35_c, x36, x38, x39, x41_c, x42, x43_c, x44_c, x45_c, x46, x49_c, x52_c, x54_c, x57, x58, x59, x61, x65, x66_c, x67_c, x70, x71_c, x72_c, x74_c, x75, x76_c, x78_c, x79_c, x80_c, x84, x85_c, x86, x88, x89_c, x90_c, x91, x93_c, x94_c, x95, x96, x98, x99_c);
and (w110, x3, x5, x6, x7_c, x19, x20, x30_c, x31, x33_c, x34, x36, x40, x43_c, x44, x47_c, x48, x54, x58, x61, x63_c, x66, x67_c, x70_c, x72_c, x76_c, x78, x81_c, x82_c, x83, x84, x89_c, x90, x93_c, x96);
and (w111, x1, x2_c, x3, x6_c, x7, x8_c, x9, x11, x12_c, x14_c, x15_c, x17_c, x18, x19_c, x20, x24_c, x27, x29_c, x31_c, x35_c, x40, x41, x42, x44, x46_c, x48_c, x49_c, x51, x52_c, x56_c, x58, x60_c, x62, x63, x68_c, x69, x71_c, x73, x74_c, x75_c, x76_c, x79_c, x81, x82_c, x84_c, x85_c, x88_c, x89_c, x93_c, x94_c, x95_c, x96_c, x97, x99_c);
and (w112, x2, x3, x4, x6, x7, x8, x9_c, x12, x14, x15, x16_c, x17_c, x18, x19_c, x20_c, x21, x22_c, x24, x25, x26, x27_c, x28_c, x29_c, x30_c, x33, x35, x36, x38, x40_c, x42_c, x44_c, x45_c, x47_c, x48_c, x49_c, x50, x51_c, x55_c, x56_c, x57_c, x58, x59, x61, x62_c, x64_c, x65, x67, x68, x69, x70, x71, x72, x73, x77, x78_c, x79, x80, x81_c, x82, x84, x86_c, x88, x89_c, x90_c, x91_c, x93, x94_c, x95, x96);
assign w113 = x89_c;
and (w114, x0_c, x1, x2_c, x3_c, x4, x6, x8, x13, x16, x17, x19, x20, x22, x24, x25_c, x26_c, x27_c, x29_c, x31, x32, x33, x34_c, x35_c, x37_c, x38_c, x39_c, x40_c, x43, x44, x45, x46_c, x47_c, x49, x52, x53_c, x54_c, x55, x56_c, x58, x61, x63_c, x64, x67, x68, x70, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x84_c, x85_c, x88, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x97, x98_c);
and (w115, x30, x36, x40_c, x55, x60_c, x63, x67, x73, x95_c);
and (w116, x0, x1, x2_c, x7, x10, x12_c, x14_c, x20, x21_c, x23_c, x24_c, x25, x26, x29, x33, x36, x37, x38, x41, x49, x54_c, x62_c, x72, x74, x76_c, x77, x80, x81_c, x83, x86_c, x87, x89_c, x94_c, x95, x96, x97, x98);
and (w117, x0_c, x1_c, x2_c, x3_c, x4_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13_c, x14, x15_c, x16, x17, x18, x19_c, x21_c, x22, x23, x25_c, x27, x28, x29_c, x30, x31, x32_c, x33, x34, x35, x36, x37_c, x38_c, x39, x41, x43, x44_c, x45_c, x46, x47, x48_c, x49, x51, x53, x54_c, x56_c, x58, x59, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69, x70, x71_c, x72_c, x73_c, x74_c, x75, x77, x78_c, x79, x81_c, x82_c, x83, x84_c, x85_c, x87_c, x89_c, x90, x91_c, x92_c, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w118, x0, x1, x3_c, x11_c, x12, x14, x19_c, x21_c, x22_c, x25_c, x27, x28, x29_c, x32_c, x33, x34_c, x35, x38, x39_c, x40, x42, x46, x47, x48_c, x50, x52_c, x54, x56, x57_c, x60, x61_c, x62_c, x63, x65_c, x66_c, x69_c, x70, x73, x76_c, x77_c, x80, x84, x88_c, x90_c, x91_c, x92_c, x93, x94_c, x97, x98);
and (w119, x1_c, x4, x13, x17, x20, x29_c, x32, x37, x60, x65, x67_c, x69_c, x75, x76_c, x84_c, x91_c, x94);
and (w120, x6, x7, x11_c, x13, x15_c, x16_c, x17, x18_c, x26_c, x29, x31_c, x33_c, x34_c, x40_c, x41, x43_c, x44, x45, x47, x49_c, x50_c, x51, x52, x58, x59, x64_c, x66_c, x67, x71, x72_c, x75_c, x78, x81_c, x83, x87, x90_c, x91, x92, x94, x95, x96, x98_c, x99_c);
and (w121, x1_c, x3, x4, x8, x9_c, x11, x13_c, x14_c, x15_c, x16, x17, x23_c, x24_c, x29_c, x30, x31_c, x35_c, x38_c, x39_c, x40, x44, x45_c, x46, x49_c, x52_c, x53, x56_c, x62, x64, x65_c, x66, x68, x72_c, x73_c, x76_c, x78, x79_c, x81_c, x83_c, x84, x86_c, x87, x88_c, x89, x90_c, x91, x92_c, x99);
and (w122, x0_c, x4_c, x7_c, x9, x14_c, x20, x22_c, x23, x24_c, x27, x30_c, x31, x36_c, x39, x40, x43, x45, x46, x47_c, x51_c, x52_c, x53_c, x57, x58, x66_c, x69_c, x70, x71, x72_c, x73_c, x78, x83, x84_c, x86, x88, x90, x93, x94, x96_c, x97, x98);
and (w123, x4_c, x7_c, x13, x18_c, x19_c, x20, x21_c, x23_c, x25, x30_c, x32_c, x37_c, x59, x67, x68_c, x73_c, x74_c, x88_c, x93, x94_c, x95);
and (w124, x0, x6_c, x7_c, x14, x16, x19_c, x22_c, x25_c, x29, x33_c, x34_c, x36, x37_c, x39, x42_c, x44, x47, x49_c, x57, x58_c, x59, x61, x62, x67_c, x70, x71_c, x72, x75_c, x78, x79_c, x83, x86, x90_c, x91_c, x95, x98_c);
and (w125, x84_c, x90_c);
and (w126, x0_c, x1, x4_c, x5_c, x6, x8, x10_c, x12, x14, x16_c, x18_c, x19, x20_c, x21, x22_c, x23_c, x25, x27_c, x29_c, x30, x33, x34, x36_c, x38_c, x39, x44, x45, x47, x49_c, x51, x52, x54_c, x56, x59, x61, x62_c, x63, x66, x67, x68, x69_c, x70_c, x75_c, x77, x78, x79_c, x80_c, x83_c, x84, x86, x87, x89, x90, x91, x92, x93_c, x94, x95, x96_c, x97, x99);
and (w127, x0_c, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x11, x12_c, x13, x14_c, x15_c, x16, x17, x18, x19_c, x20_c, x22_c, x23_c, x24_c, x25_c, x26_c, x28, x29_c, x30, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37, x38_c, x39, x40, x41_c, x42_c, x43, x44, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x54, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63, x64_c, x65, x68_c, x69, x70_c, x73, x74, x75, x76, x77, x78_c, x79_c, x80, x81_c, x82, x83, x85_c, x86, x87, x88, x89_c, x90_c, x91, x92_c, x94, x95, x96_c, x97, x98, x99);
and (w128, x0_c, x2, x3_c, x6, x7, x8_c, x11_c, x12, x14, x15_c, x17, x22, x25_c, x26_c, x27, x32_c, x39_c, x42, x48_c, x50, x56_c, x64_c, x65_c, x67_c, x78, x80, x83, x84_c, x85_c, x86, x89, x90_c, x92_c, x94_c);
and (w129, x1_c, x2, x3_c, x4, x5_c, x6_c, x8_c, x9_c, x10_c, x11_c, x14, x16_c, x18, x20, x22_c, x23, x24, x25, x28_c, x30_c, x31, x32_c, x33, x37, x39, x40, x41_c, x43, x45_c, x46_c, x47, x49, x50, x51, x52, x53, x55, x56, x57_c, x58_c, x59_c, x60, x62, x63_c, x64_c, x66_c, x67, x68_c, x70_c, x71, x72, x74, x75_c, x77, x78, x80, x81, x82, x83, x84, x85, x86_c, x87_c, x89, x90_c, x91, x93_c, x94_c, x95, x97_c);
and (w130, x1_c, x4, x8, x33_c, x44_c, x69, x81, x85, x91, x97_c);
and (w131, x2_c, x3_c, x4, x5_c, x6_c, x7, x8_c, x9_c, x11_c, x12_c, x13, x15_c, x16_c, x17, x18, x19, x20, x22, x23, x24_c, x25, x27, x29, x30, x31_c, x34, x35, x36_c, x37, x39, x40, x41, x42, x43_c, x44, x45_c, x46, x48_c, x49_c, x50, x51_c, x52, x54, x55, x57, x58, x59_c, x61, x62, x65, x66, x67_c, x68, x69, x70, x72, x73_c, x74, x75_c, x77_c, x79_c, x80, x81, x82_c, x83, x84, x86, x88_c, x90, x91, x92, x93_c, x94_c, x95, x98, x99);
and (w132, x0_c, x1_c, x2, x3_c, x8_c, x10, x11_c, x12, x16, x18_c, x20, x21, x22, x23, x26, x27, x30, x31, x32_c, x33, x34, x39_c, x44_c, x47, x55_c, x58, x60, x62, x66_c, x67, x69_c, x74, x75_c, x77_c, x82_c, x85, x93_c, x95_c, x98, x99_c);
and (w133, x0, x1_c, x2_c, x4, x5_c, x6, x8_c, x10_c, x13, x14_c, x17_c, x18, x19, x20, x24, x25_c, x27_c, x28_c, x29, x30_c, x33_c, x34_c, x36, x37, x38, x40, x41_c, x46_c, x47, x49_c, x50_c, x52_c, x53, x54_c, x55_c, x56, x57_c, x63_c, x64, x65_c, x66, x67, x68, x70, x71, x73_c, x74_c, x75, x76_c, x77, x78_c, x79_c, x80_c, x83_c, x84, x85, x88, x89_c, x91_c, x92, x94, x95_c, x96, x97_c, x98_c, x99);
and (w134, x0, x1, x2, x3, x4, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13, x14_c, x16, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26_c, x27, x28_c, x29, x30, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48_c, x49_c, x50, x51_c, x52, x53, x54_c, x55_c, x56, x57_c, x58, x59_c, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x67, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80, x81_c, x82_c, x83, x84_c, x85, x86, x87_c, x88, x89, x90, x91_c, x92_c, x94_c, x95, x96_c, x97, x98, x99);
and (w135, x1_c, x2, x5_c, x6, x11_c, x12, x14, x15, x19_c, x26_c, x27, x30, x32_c, x35, x39, x41_c, x42_c, x43, x49, x55, x62_c, x63, x64_c, x67_c, x70_c, x71_c, x72, x75, x76, x79, x80_c, x82, x84, x85_c, x89, x90_c, x93, x96);
and (w136, x1_c, x3, x10_c, x11, x12, x15_c, x16_c, x18_c, x20_c, x22, x23_c, x24, x26, x28_c, x29, x35, x36, x39_c, x41, x43_c, x45_c, x46, x48, x49_c, x51, x52_c, x53_c, x56_c, x57_c, x60_c, x61, x64, x67, x68_c, x69_c, x73, x74, x75, x79, x81_c, x85, x86, x90_c, x92_c, x96, x97, x99_c);
and (w137, x0_c, x1, x3_c, x5_c, x6, x7, x9_c, x10_c, x11, x12_c, x14, x16_c, x17_c, x22_c, x23, x26_c, x28_c, x29, x32_c, x33, x35_c, x36_c, x38, x39_c, x40_c, x41_c, x43, x44, x46_c, x49_c, x50, x54, x55_c, x57, x64_c, x67_c, x71_c, x73, x74, x75_c, x76, x78, x79, x81_c, x82, x84, x86, x87_c, x89_c, x91, x93_c, x96, x99_c);
and (w138, x1, x3, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x12, x13, x14_c, x15, x16, x17_c, x18, x19, x20_c, x22_c, x23_c, x24_c, x25, x26, x27_c, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35, x36, x38, x39, x41, x42, x43_c, x44, x45_c, x46_c, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55_c, x56, x58_c, x60, x61_c, x62, x63, x64_c, x65, x66_c, x68, x69, x70_c, x71_c, x72, x73_c, x74_c, x75, x76, x78, x79_c, x80, x81_c, x82_c, x84, x85_c, x86_c, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94_c, x96, x98_c, x99_c);
and (w139, x1, x7, x8_c, x10, x17_c, x23, x26_c, x34, x40, x46, x48_c, x49_c, x58_c, x61_c, x62, x68_c, x69, x72, x74, x80_c);
and (w140, x0, x2_c, x3_c, x5, x6, x8, x10_c, x11_c, x13_c, x14, x15, x17_c, x18, x20_c, x23, x24, x25, x27, x28_c, x29, x31_c, x34_c, x35_c, x36, x38_c, x39, x43, x45_c, x48, x49_c, x51_c, x52_c, x54_c, x55, x56_c, x57_c, x60, x61, x62, x63, x65_c, x67, x70, x71_c, x72_c, x73, x74, x76_c, x78, x82, x85, x88, x90, x91_c, x92_c, x93_c, x96_c, x97, x98_c, x99);
and (w141, x39_c, x54, x55, x58_c, x62, x71, x81_c, x94);
and (w142, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14, x15_c, x16, x17_c, x18, x19_c, x20, x21_c, x22, x23, x24, x25_c, x26, x27, x28_c, x29, x30, x31_c, x32, x33_c, x34_c, x35, x36_c, x37_c, x38_c, x39_c, x40, x41, x42_c, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56, x57, x58, x59_c, x60_c, x61_c, x62, x63, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x81, x82_c, x83, x84, x85, x86_c, x87, x88_c, x89, x90_c, x91, x92, x93, x94, x95, x96_c, x97_c, x98, x99);
and (w143, x0, x2, x3_c, x4_c, x5, x6, x7, x8, x9_c, x10_c, x11, x12, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20, x21_c, x23, x24, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38_c, x39, x40, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47, x48, x49, x50_c, x51, x52_c, x53, x54, x55_c, x56_c, x57, x58, x59_c, x60, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68, x69, x70_c, x71, x72, x73_c, x74_c, x75, x76, x77_c, x78, x80, x81, x82_c, x83_c, x84_c, x85_c, x86, x87, x88_c, x90, x91_c, x92, x93, x94, x95, x96, x97, x98);
and (w144, x2_c, x4, x5, x7_c, x9_c, x13_c, x14_c, x18_c, x19, x20_c, x22_c, x24_c, x28_c, x30, x32, x35_c, x36_c, x37_c, x38, x40, x44, x47_c, x48, x50, x52_c, x59, x61_c, x63_c, x65, x71_c, x72, x73, x76_c, x77, x79_c, x80, x81, x83, x84, x87_c, x89_c, x93, x94_c, x97, x98);
and (w145, x1_c, x2_c, x4, x7_c, x8, x9, x11, x15, x16_c, x19, x22_c, x26, x28, x30, x31_c, x32_c, x35_c, x39_c, x44, x45, x46, x57, x58, x61_c, x62_c, x65_c, x66, x67, x68_c, x70, x71_c, x73_c, x75_c, x76_c, x78, x81, x82_c, x83_c, x84, x85_c, x87, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95_c, x99_c);
and (w146, x4_c, x20_c, x25_c, x33_c, x34, x41_c, x43_c, x46_c, x50, x54, x66, x69, x72_c, x77_c, x80, x82, x86);
and (w147, x2_c, x21, x62, x81_c, x98);
and (w148, x7, x22, x29, x36, x37_c, x40_c, x41_c, x44, x47, x48_c, x49_c, x53, x56_c, x67_c, x68_c, x78_c, x79, x84, x89_c, x90_c);
and (w149, x1_c, x3_c, x4, x5, x7_c, x8, x9, x11_c, x13_c, x14, x16_c, x17, x18, x20, x21, x22_c, x26_c, x27_c, x28, x35, x38_c, x39, x41_c, x52_c, x57, x59_c, x72_c, x74_c, x77_c, x78, x80, x85_c, x88, x93_c, x98);
and (w150, x0, x1, x2_c, x3, x5, x6, x7, x8, x9_c, x11, x12, x13_c, x14_c, x15, x16, x17_c, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x24, x26, x28_c, x29, x30, x31, x32_c, x34, x36, x40, x41_c, x42, x46_c, x47, x49_c, x50, x52_c, x53_c, x54, x55_c, x56_c, x58, x60, x64, x65_c, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73_c, x74, x76, x78, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91_c, x92_c, x93, x94, x95_c, x96, x98, x99_c);
and (w151, x0_c, x3_c, x6, x7, x8_c, x9_c, x12_c, x13_c, x14_c, x15, x16, x19, x20_c, x21_c, x22_c, x24, x25, x26_c, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x38_c, x39, x41, x42_c, x43, x45, x46_c, x47, x48, x49_c, x50, x51, x52_c, x53, x54, x55_c, x57_c, x58_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x67, x68_c, x70, x71_c, x72, x75, x76, x77_c, x78, x79_c, x80_c, x85_c, x87, x89, x91_c, x92, x93, x94, x95_c, x96, x97, x98, x99);
and (w152, x14_c, x28, x30_c, x31, x35, x42, x46_c, x53, x54, x55, x76_c);
and (w153, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10_c, x12_c, x14, x16, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34_c, x38_c, x39_c, x40, x41_c, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x53_c, x55_c, x56, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69_c, x70, x72, x73_c, x74_c, x76, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85, x86, x87, x88_c, x91, x92, x93_c, x94_c, x95, x96, x97, x98_c, x99_c);
and (w154, x14, x15, x20_c, x31_c, x36_c, x42_c, x48, x59_c, x63, x64, x67_c, x70, x73_c, x74_c, x88);
and (w155, x1_c, x4_c, x7_c, x9, x10, x13_c, x14_c, x15_c, x16, x17_c, x20, x25_c, x28_c, x29, x30_c, x31_c, x32_c, x34, x35_c, x36_c, x37_c, x39, x43, x47, x49_c, x52_c, x53_c, x54_c, x56, x65_c, x66, x68_c, x70_c, x73_c, x74, x78_c, x80, x84, x89, x90, x93_c, x99);
and (w156, x0, x1, x3, x4, x5, x6_c, x7, x8, x9, x10, x11_c, x12_c, x13_c, x14_c, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23_c, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32_c, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40, x41, x42_c, x43, x44, x45_c, x46, x47, x48, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57, x58, x59, x60, x61_c, x62, x63, x64, x65_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85, x86_c, x87, x88, x89_c, x90, x91, x92_c, x93, x94, x95_c, x96, x97_c, x98, x99_c);
and (w157, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8_c, x10_c, x12, x13, x14, x15_c, x16_c, x17_c, x18_c, x19, x20_c, x21, x22, x23_c, x24, x25, x26_c, x27_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36_c, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49_c, x50, x51_c, x52, x53, x54, x55, x56, x57, x58_c, x59, x60, x61_c, x63, x64_c, x66_c, x68, x69, x70_c, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x79, x81_c, x82, x84, x85, x86, x87, x88, x89_c, x90_c, x91, x92_c, x93, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w158, x13_c, x49, x64, x71, x72_c, x79);
and (w159, x1_c, x4, x5_c, x6_c, x7_c, x10_c, x14_c, x16, x17_c, x19_c, x20, x22_c, x25, x26_c, x27_c, x28, x30_c, x32, x33, x34_c, x35_c, x37, x38_c, x41, x43_c, x44, x48_c, x51, x52, x53, x55, x56, x58, x59_c, x60_c, x66, x70, x71_c, x73, x78_c, x79_c, x81_c, x82_c, x83, x84, x86, x88, x89, x92, x93_c, x94_c, x96_c, x97_c, x99);
and (w160, x9, x10, x16_c, x17_c, x21_c, x25_c, x38_c, x55, x61_c, x63, x83, x89, x96);
and (w161, x21_c, x35_c, x41, x57, x59_c, x62_c, x73_c, x85_c, x91);
and (w162, x0, x1, x3, x4_c, x5_c, x7, x8, x9, x12_c, x13, x14_c, x15, x17_c, x18, x19_c, x20, x22, x23, x24_c, x25, x26_c, x28_c, x29, x30, x33, x34, x35, x36_c, x37, x38_c, x39, x40, x42_c, x43, x45_c, x47, x48, x51, x52, x53, x55_c, x56_c, x57, x58, x59_c, x61_c, x65_c, x66_c, x67_c, x68_c, x72, x73_c, x74, x76, x77_c, x78, x81, x82, x83, x84_c, x85, x88, x90, x91_c, x92, x93_c, x95_c, x96_c, x97, x98, x99_c);
and (w163, x2_c, x3_c, x11, x17, x20_c, x25_c, x27_c, x30, x39_c, x42, x43, x50_c, x53_c, x74, x79, x87_c, x91, x93);
and (w164, x0_c, x1, x9, x10_c, x20, x23, x31_c, x35, x39_c, x42_c, x44_c, x47, x50_c, x62, x65_c, x73_c, x76, x77, x79, x81, x83_c, x84_c, x87_c, x91, x99);
and (w165, x1, x3_c, x7_c, x9, x12_c, x13_c, x14, x16, x19, x20, x23, x25, x27, x28, x31, x33_c, x35_c, x39_c, x40_c, x41, x43_c, x47, x48_c, x49_c, x50_c, x52_c, x54, x55, x56, x58, x59_c, x66, x69, x73_c, x74_c, x76, x77, x81_c, x82_c, x83_c, x86, x87_c, x88, x89, x91_c, x92, x95_c);
and (w166, x0_c, x1_c, x2_c, x3_c, x4, x5, x6, x7_c, x8_c, x9_c, x10_c, x12_c, x13, x14_c, x15, x16_c, x17, x18_c, x19_c, x20, x22_c, x23, x24_c, x25, x26, x27_c, x28_c, x29_c, x30, x31, x32_c, x33_c, x34_c, x36, x38_c, x39, x40_c, x41, x42_c, x43, x44, x45_c, x46, x47, x48_c, x50, x51, x52, x53_c, x54_c, x55, x56, x57, x58, x59, x60, x61_c, x62, x64_c, x65_c, x66_c, x67, x69_c, x70_c, x71_c, x72_c, x73, x74_c, x75_c, x76_c, x77_c, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87_c, x88, x89, x90, x91, x92_c, x93_c, x94_c, x95_c, x96_c, x97, x98, x99);
and (w167, x2, x4, x18_c, x26_c, x30_c, x33, x39, x55_c, x57, x59_c, x66_c, x72_c, x74_c, x88, x92, x94_c, x95, x99);
and (w168, x0, x1, x2, x3_c, x4, x5, x6, x7_c, x8_c, x9, x10, x12, x13, x14, x15, x17_c, x18, x19, x20_c, x21, x24_c, x25_c, x26_c, x27_c, x32, x33_c, x34_c, x35, x36, x38, x40_c, x42_c, x45_c, x46, x47, x49_c, x50_c, x51_c, x54_c, x59_c, x60, x61, x63, x64, x65, x66_c, x68_c, x70_c, x71_c, x72_c, x73_c, x74, x76, x77_c, x78, x79_c, x80, x83, x87_c, x88_c, x89_c, x90, x92, x94_c, x97_c, x99_c);
and (w169, x1_c, x2, x4_c, x6_c, x10, x13_c, x14_c, x19_c, x20, x21_c, x23, x24_c, x28_c, x29, x31, x34_c, x35_c, x36_c, x40_c, x42, x47_c, x48_c, x49, x50, x51_c, x53_c, x54, x55, x57_c, x58_c, x61_c, x62_c, x63_c, x65, x66_c, x67, x69_c, x70, x71, x73, x75, x76_c, x77, x80, x82_c, x83_c, x84, x85_c, x86, x89, x95);
and (w170, x0, x2, x6, x7, x8, x9_c, x10, x13_c, x15_c, x16_c, x18_c, x19, x20_c, x22, x25_c, x27, x29, x30, x31_c, x32_c, x34_c, x35_c, x37, x41_c, x42_c, x43_c, x44, x45_c, x46_c, x47, x49, x54_c, x55, x56, x57_c, x62_c, x63, x66, x68, x74_c, x80, x81_c, x82_c, x84, x88_c, x89, x91, x94_c, x99_c);
and (w171, x0, x1, x6_c, x7, x10_c, x12_c, x14_c, x15, x17_c, x18_c, x21, x24_c, x25, x28, x30, x32, x36_c, x39, x41_c, x44, x48, x51_c, x54, x55, x56, x58_c, x59, x60_c, x61, x62, x64_c, x65, x66_c, x68_c, x69_c, x70, x73_c, x74, x77, x79, x81_c, x82, x83, x87, x88, x89_c, x92_c, x93_c, x94, x95_c, x97_c, x98, x99);
and (w172, x0, x2, x3_c, x4, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16_c, x17_c, x18, x19, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x28_c, x29_c, x30, x31_c, x32, x33_c, x34_c, x35, x36_c, x37_c, x38, x39_c, x40, x41, x42, x43_c, x44, x45_c, x46, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58_c, x60, x61_c, x62_c, x63, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80, x81_c, x82, x83_c, x84_c, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91_c, x92, x93, x94_c, x96_c, x97, x98_c, x99);
and (w173, x5, x6, x7_c, x10, x11_c, x13, x20_c, x24, x29, x32_c, x37_c, x39_c, x40, x41_c, x44, x45, x46_c, x47, x52_c, x59_c, x60_c, x61_c, x63_c, x66_c, x67, x70, x72, x79, x81_c, x84_c, x85, x88, x89, x91, x96, x99_c);
and (w174, x0, x1, x2_c, x3_c, x6_c, x7_c, x9, x11, x12, x14, x16, x17_c, x18_c, x19_c, x20, x21_c, x22, x23, x24, x25_c, x26, x27_c, x28, x29, x30, x31_c, x32, x33, x34_c, x35_c, x36_c, x37, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52_c, x53, x54, x56_c, x57, x58_c, x59, x60, x61_c, x62, x63_c, x64, x65, x66, x67, x68, x69, x70_c, x71_c, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x84, x85, x86, x88, x89_c, x90_c, x91_c, x94, x96, x97_c, x98_c, x99_c);
and (w175, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x7, x9_c, x10_c, x14, x16_c, x18, x19_c, x20, x21, x23, x24, x25_c, x26_c, x27, x28_c, x29, x30, x31_c, x32, x33_c, x34_c, x35, x36, x37_c, x38_c, x40, x41_c, x44_c, x45, x46_c, x50_c, x51, x52_c, x53_c, x54, x55_c, x56_c, x57, x58, x59, x61, x62, x63, x64_c, x66, x67, x68, x69, x71_c, x72_c, x73, x75_c, x77, x79, x80_c, x81, x82, x83, x84, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93, x98_c);
and (w176, x0_c, x1, x3, x5, x6, x7, x9, x10_c, x13, x15_c, x17_c, x21_c, x24_c, x26_c, x28, x30, x31, x33_c, x36_c, x41, x45_c, x46_c, x47_c, x54, x56, x61_c, x64, x66_c, x67_c, x75, x78_c, x85, x86, x87_c, x88, x89_c, x94_c, x96, x97_c);
and (w177, x0, x2, x3, x4, x7, x10, x13_c, x14_c, x17_c, x19, x20, x21, x24, x25, x27_c, x28_c, x29, x30_c, x31_c, x32_c, x33_c, x35_c, x36_c, x40, x41, x42_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x52_c, x54, x56, x57_c, x58, x59_c, x60_c, x62_c, x64_c, x65_c, x66, x67, x69_c, x70_c, x72_c, x73, x74, x75, x77_c, x78_c, x79_c, x80, x81, x82, x83_c, x84_c, x85_c, x86, x87_c, x88_c, x89_c, x91_c, x92, x93_c, x94, x95_c, x96, x97_c, x98, x99);
and (w178, x3, x4, x5_c, x6, x7, x8, x10_c, x14_c, x16_c, x17, x18, x24_c, x25_c, x27, x28, x29, x31, x34, x36, x37, x38_c, x41_c, x42_c, x45, x47, x48, x49, x53_c, x54, x57_c, x58_c, x59_c, x60_c, x63_c, x64_c, x66_c, x67_c, x68_c, x69, x74_c, x76_c, x78, x81, x82_c, x85_c, x91_c, x92, x96_c, x98_c, x99_c);
and (w179, x8, x32_c, x57, x76_c, x79_c, x97_c);
assign w180 = x13_c;
and (w181, x0_c, x2_c, x3_c, x5_c, x6_c, x8, x9_c, x10, x11_c, x12, x13_c, x14, x15_c, x16_c, x18, x19, x20_c, x21_c, x22, x23, x24, x25, x26_c, x27_c, x28_c, x29_c, x30, x31_c, x32, x33_c, x34, x35, x36, x37, x38_c, x39, x41_c, x42_c, x43, x44, x45_c, x47, x48_c, x49, x50_c, x51, x53, x54_c, x55_c, x57_c, x58, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66, x67, x69_c, x70_c, x71, x73_c, x74, x75, x76, x79, x80_c, x82_c, x83, x84, x85, x88_c, x89_c, x90, x91_c, x93, x95_c, x96_c, x97, x98, x99_c);
and (w182, x0, x1, x2_c, x3, x4_c, x5, x6, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15, x16, x17, x18, x19, x20, x21, x22_c, x23_c, x24, x25, x26_c, x27_c, x28, x29_c, x30_c, x31_c, x32, x33, x34, x35_c, x36, x37_c, x38_c, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x51, x52_c, x53, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61, x62_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69, x70, x71_c, x72, x73_c, x74_c, x75, x76, x77_c, x78, x79_c, x80, x81_c, x82, x83_c, x85, x86_c, x87_c, x88_c, x89, x90, x91, x92_c, x93_c, x94_c, x95_c, x96, x97, x98_c, x99_c);
and (w183, x0, x1, x2, x3, x4, x5_c, x7_c, x8_c, x9_c, x10_c, x13, x14, x15_c, x16, x17, x18, x19_c, x23, x24, x25, x26_c, x27, x28, x29, x30, x31_c, x32_c, x33, x34_c, x36_c, x37, x39, x43_c, x44, x45_c, x46_c, x47, x48, x50_c, x51, x52, x53_c, x54_c, x55_c, x56_c, x58, x59_c, x62, x63_c, x64, x65, x67, x69_c, x70, x71_c, x73_c, x74, x75_c, x76, x79, x80_c, x81, x82, x84, x85, x86_c, x87_c, x92, x93, x94_c, x95, x97_c, x98, x99_c);
and (w184, x0, x2_c, x3, x4_c, x5_c, x7_c, x9_c, x12_c, x13, x14, x15, x17_c, x18, x19_c, x20, x21, x22, x23, x25, x28_c, x29_c, x31, x32_c, x35, x39_c, x40_c, x41, x42, x43, x45, x47_c, x49, x51, x52_c, x54, x55_c, x56_c, x59_c, x60, x62, x63, x64, x65, x66_c, x67_c, x68_c, x69, x71_c, x73_c, x74_c, x75, x76_c, x78_c, x79, x80, x81_c, x84_c, x86, x87_c, x89, x90_c, x92_c, x93, x96_c, x98_c, x99_c);
and (w185, x3_c, x6, x7, x22_c, x25_c, x28_c, x32, x35, x37, x40, x45_c, x46, x47_c, x50, x56, x63_c, x66_c, x67_c, x69, x71, x75, x81_c, x84, x92_c);
and (w186, x0, x3, x53_c, x59_c, x77, x82_c, x91);
and (w187, x1_c, x2, x6_c, x8_c, x14, x17, x21, x22, x28, x32, x33_c, x36, x41, x43_c, x44_c, x46_c, x49, x63_c, x65, x72, x73, x75, x76_c, x87_c, x91_c, x97_c, x99_c);
and (w188, x4, x5_c, x6, x8_c, x11_c, x12, x13_c, x14_c, x15_c, x17_c, x19_c, x20_c, x27_c, x30_c, x31, x32, x35, x36, x37_c, x39_c, x40, x42, x50_c, x54, x56_c, x58, x63, x65, x69, x70, x71_c, x73_c, x74, x76_c, x77_c, x78_c, x79, x83, x87_c, x90, x91_c, x95, x96, x97, x99_c);
and (w189, x0_c, x1_c, x2_c, x3, x4, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16_c, x17, x19_c, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x33_c, x34, x36, x37_c, x38, x39, x40, x41, x43_c, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81, x82, x83, x85_c, x86_c, x87, x88_c, x89, x90, x92, x94, x95, x97_c, x98, x99_c);
and (w190, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7, x8, x9_c, x10_c, x11, x12, x13_c, x14_c, x15, x16_c, x17_c, x18, x20_c, x21_c, x22_c, x23_c, x25_c, x26, x27_c, x28, x29, x30_c, x31_c, x32, x33, x34_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x41, x42, x43_c, x44_c, x45, x46_c, x47_c, x48, x49, x51, x52, x53, x54_c, x55, x56_c, x57_c, x58, x59_c, x60_c, x61_c, x62, x64_c, x65_c, x66_c, x67_c, x68, x69, x70, x71_c, x72, x73_c, x74, x75, x76_c, x77, x78_c, x79_c, x80_c, x81_c, x82, x83, x84, x85, x86_c, x87, x88, x89, x90_c, x91, x92_c, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w191, x0, x2, x3_c, x5, x6_c, x9_c, x12, x13, x14_c, x16_c, x18, x21_c, x24_c, x25, x31_c, x35_c, x37, x40, x41_c, x43, x44_c, x45_c, x46, x47_c, x48, x49_c, x51_c, x52, x54, x55_c, x57_c, x58, x59, x60_c, x63_c, x64, x65, x67, x69_c, x72, x73, x75_c, x77, x78, x80, x82, x84, x88_c, x89_c, x92_c, x93_c, x94, x97, x98, x99);
and (w192, x1_c, x2, x3_c, x4, x7_c, x9, x11_c, x12_c, x14_c, x15, x19, x20, x22, x24_c, x25_c, x28_c, x31, x32_c, x36, x37_c, x38, x42, x46, x48, x49_c, x52, x54_c, x56_c, x64, x68, x73_c, x76, x77, x79, x81_c, x83, x85, x86, x88, x90_c, x91);
and (w193, x0, x4, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x12, x13, x14, x16_c, x17, x19_c, x20, x21_c, x22_c, x23, x24, x26_c, x27, x29_c, x30, x31_c, x33_c, x34_c, x35, x36_c, x37_c, x38, x39_c, x40, x41, x43_c, x44, x46, x48, x49, x50, x51, x52, x53_c, x54_c, x55, x56, x57, x58, x60_c, x63, x64_c, x65, x66_c, x67_c, x68, x70, x71, x72, x73, x74, x75_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84, x88, x89_c, x90_c, x91_c, x92, x94, x95_c, x96_c, x97, x99_c);
and (w194, x0, x6, x9, x11_c, x14, x15_c, x21, x22, x24, x31, x33_c, x35_c, x41, x44_c, x49, x53, x60, x62, x65_c, x66_c, x79, x83, x91_c, x93_c, x94_c);
and (w195, x0_c, x2, x3_c, x5, x7, x9_c, x11, x13, x16_c, x19_c, x22, x23_c, x24_c, x27_c, x28_c, x31_c, x32, x36_c, x38, x43, x49_c, x50_c, x52_c, x53, x56_c, x58, x59_c, x62_c, x64, x65, x66_c, x67_c, x68_c, x72_c, x73, x78, x83, x84_c, x88, x91, x93, x96, x97, x98_c, x99_c);
and (w196, x0_c, x1, x2_c, x3_c, x4, x5, x6_c, x7, x8, x9, x10_c, x11_c, x12_c, x13, x14_c, x15_c, x16, x17_c, x18_c, x19, x20, x21_c, x22_c, x23_c, x24, x25, x26_c, x27, x28_c, x30_c, x31, x32_c, x33_c, x34_c, x36_c, x37_c, x39_c, x40, x41_c, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50_c, x51, x52_c, x53, x54, x55_c, x56_c, x57_c, x58, x60, x61, x62_c, x63, x64, x65_c, x66, x67, x68_c, x69, x70, x71_c, x72, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84, x85_c, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94_c, x95_c, x96_c, x97, x98, x99_c);
and (w197, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x23_c, x25_c, x27_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x47_c, x48, x53, x54_c, x56_c, x58_c, x59_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80_c, x82, x84_c, x85, x86, x87_c, x89, x90, x91_c, x92, x93_c, x96, x98_c, x99);
and (w198, x0, x1_c, x2_c, x3, x4_c, x6_c, x7_c, x8, x10, x11_c, x12_c, x13, x14, x15, x16, x17_c, x20_c, x22, x23_c, x25_c, x26_c, x27, x28, x29, x30_c, x31_c, x33_c, x34, x36, x37_c, x39_c, x40_c, x42_c, x43, x46, x47_c, x48_c, x49, x50, x51_c, x52_c, x53, x54, x55_c, x56, x57_c, x58_c, x59, x61_c, x62, x63_c, x64, x65_c, x68_c, x69_c, x71_c, x72_c, x73, x74_c, x75_c, x77, x78_c, x79_c, x82_c, x83_c, x84_c, x85, x87, x88_c, x89, x91_c, x92_c, x93, x94, x95, x96_c, x97_c, x98, x99_c);
and (w199, x0_c, x1_c, x5, x8, x10, x11_c, x20_c, x23, x30, x33_c, x35, x36_c, x37_c, x47_c, x48, x60_c, x62_c, x64_c, x69_c, x70, x72_c, x73, x77, x78_c, x79_c, x83_c, x85_c, x86, x90_c, x92);
and (w200, x0_c, x2_c, x5_c, x7_c, x8_c, x9, x10, x11_c, x13_c, x14_c, x20, x21_c, x23, x24, x25_c, x26, x27, x28_c, x29_c, x30, x32, x33, x36, x37, x38, x39, x40, x45_c, x49, x50, x53_c, x54_c, x55_c, x57, x58_c, x60_c, x61, x62_c, x63_c, x64, x72_c, x73_c, x77_c, x78_c, x80_c, x81_c, x84, x86, x87_c, x91, x92, x93_c, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w201, x26, x33_c, x44, x53);
and (w202, x2_c, x19, x24_c, x26, x36, x46_c, x55_c, x92_c, x95_c, x98);
and (w203, x0_c, x1, x2, x3_c, x4_c, x5_c, x7_c, x8, x10_c, x11_c, x12_c, x13, x14_c, x16_c, x17_c, x18_c, x20_c, x21, x22_c, x24, x26, x27_c, x28_c, x29_c, x30, x31_c, x32_c, x34, x35_c, x36_c, x39_c, x40, x41, x42_c, x43, x44, x46, x47, x48_c, x49_c, x50, x51_c, x53_c, x54_c, x56_c, x57, x58, x59, x60_c, x62, x63_c, x65, x66_c, x67, x68_c, x69, x70, x71, x73_c, x74, x75, x76, x77_c, x78, x79, x80, x81_c, x82, x85_c, x88, x90_c, x91, x93, x95, x96, x97_c, x98_c);
and (w204, x0, x2_c, x3, x4_c, x5_c, x6_c, x7, x10_c, x11, x12, x13, x14, x17, x18_c, x20_c, x21_c, x22_c, x24, x25_c, x26_c, x27, x28_c, x31_c, x32, x34, x35, x38, x39, x41, x44_c, x45_c, x46, x47, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58, x59, x60_c, x61, x62, x63, x64_c, x65_c, x66_c, x67, x68_c, x69, x71_c, x73, x75, x77, x78, x79_c, x80, x81, x83_c, x84_c, x85_c, x86_c, x88, x90_c, x91_c, x92_c, x93_c, x95, x98_c);
and (w205, x0, x2, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x11_c, x12_c, x13, x14_c, x15_c, x16, x17_c, x18, x19_c, x20_c, x21, x22, x26, x27_c, x28, x29, x30, x31, x32, x34, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41, x42_c, x44, x45, x46_c, x47, x48, x49, x51_c, x52_c, x53, x55_c, x56, x58, x59, x61_c, x63, x65, x66_c, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74, x75, x76, x77_c, x78, x79_c, x80, x81, x82_c, x83, x85_c, x86, x87_c, x89_c, x92, x93, x94_c, x95_c, x96_c, x97, x98_c, x99_c);
and (w206, x1, x3_c, x4_c, x5_c, x6_c, x7_c, x8, x9, x10_c, x11, x12, x13, x14, x15, x16_c, x18, x19, x21, x22, x23, x24_c, x26_c, x27_c, x29, x30_c, x31_c, x32_c, x33, x34, x35_c, x36_c, x37, x38_c, x40, x41, x42, x43_c, x44_c, x45, x46_c, x48, x49_c, x50_c, x52, x53, x54, x55, x56_c, x57_c, x58_c, x59, x60, x61, x62, x63_c, x65_c, x66_c, x67_c, x68_c, x70_c, x71, x72, x73, x75_c, x76, x77_c, x78, x79, x80_c, x81, x82_c, x83, x84_c, x86, x87, x88, x90, x91, x93_c, x94, x95, x96, x97, x98_c);
and (w207, x0_c, x1, x2, x3_c, x4_c, x5, x6_c, x8_c, x9, x11_c, x12, x13, x16_c, x18, x19, x20_c, x21, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29_c, x30, x31, x32, x33, x34, x35, x36, x37_c, x38_c, x39, x40, x41, x43_c, x44_c, x45_c, x46_c, x47_c, x48, x49, x50_c, x51, x52_c, x53, x54_c, x56, x57, x58_c, x59_c, x60, x62_c, x63_c, x65, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x83, x84_c, x85_c, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92, x93, x94, x95, x96_c, x97_c, x99);
and (w208, x0, x2_c, x3, x8_c, x9, x14_c, x17_c, x18, x29_c, x32, x35, x37, x38_c, x42_c, x49, x51, x52, x57, x58_c, x59, x60_c, x68, x69, x71, x75_c, x76, x78_c, x80, x89, x90_c, x98);
and (w209, x2_c, x4_c, x6_c, x7_c, x9, x11, x12_c, x14, x16_c, x18, x20_c, x21_c, x22_c, x23_c, x24, x25, x26, x27_c, x28, x32_c, x33, x36, x37_c, x39, x41, x43, x45_c, x51, x52, x53, x54_c, x56_c, x57_c, x58_c, x61, x62, x66_c, x68_c, x69_c, x71_c, x73_c, x74_c, x75, x76, x77, x80_c, x81_c, x84, x85, x86_c, x94, x96_c, x98_c, x99_c);
and (w210, x7, x16_c, x21, x24, x26, x37_c, x40, x41_c, x44, x48_c, x53, x64_c, x74, x76_c, x78_c, x80, x82_c, x86_c, x90_c, x91, x94_c, x95);
and (w211, x8_c, x49_c, x75, x89_c);
and (w212, x0_c, x2_c, x4, x6_c, x9_c, x10_c, x11, x14_c, x15_c, x16, x21, x23, x25_c, x26_c, x27, x28_c, x29_c, x31, x32_c, x33_c, x36_c, x37, x38, x41_c, x42, x43_c, x44, x45, x46, x49, x50_c, x53_c, x54, x55, x57, x59, x60_c, x65, x69_c, x72_c, x73_c, x79_c, x80, x81_c, x83, x84, x87, x89, x92_c, x93, x94, x95, x96_c, x97_c);
and (w213, x0, x2_c, x3_c, x4_c, x5, x7_c, x9, x11_c, x12, x14_c, x15_c, x18, x21_c, x22, x28, x30_c, x31, x32, x34, x35_c, x37, x38, x39_c, x43, x47_c, x49_c, x50, x51_c, x52, x55_c, x59, x60, x63, x66, x68_c, x72_c, x75_c, x76_c, x78, x82_c, x84_c, x88_c, x89, x90_c, x91, x92, x93_c, x95_c, x96);
and (w214, x0_c, x3_c, x6, x7, x10_c, x11_c, x12, x13, x15, x16_c, x18_c, x19_c, x23_c, x26, x34, x39, x40, x47_c, x49, x53, x54, x57_c, x61, x62_c, x63, x64_c, x66, x67, x69_c, x77, x78_c, x80_c, x81, x86, x87, x89_c, x90_c, x92, x94, x95, x98, x99);
and (w215, x49, x94_c, x96_c);
and (w216, x1_c, x2, x4_c, x7, x9_c, x10, x11_c, x12_c, x15, x17_c, x18, x19_c, x20, x22, x24_c, x25, x26_c, x27, x28_c, x29, x30, x31, x32, x34_c, x36_c, x39_c, x40_c, x44, x46_c, x47, x49_c, x50_c, x51, x52_c, x53_c, x55_c, x56, x58_c, x59, x60, x63, x65_c, x67_c, x68_c, x69, x70, x71, x73_c, x74, x78_c, x79_c, x80, x86, x87, x88, x89, x90_c, x93, x94, x96, x97, x98_c, x99);
and (w217, x0_c, x1, x2, x3_c, x4_c, x5, x6_c, x7_c, x8, x9_c, x11_c, x13, x14_c, x15, x17, x18, x19_c, x25_c, x26_c, x27_c, x28_c, x29_c, x30, x31_c, x32_c, x33_c, x35, x37_c, x38_c, x39, x40, x41, x42, x43_c, x44_c, x45, x47_c, x48, x49_c, x51_c, x52, x53_c, x54_c, x56_c, x57, x58_c, x59_c, x60_c, x61, x63_c, x64, x67, x68, x69, x70, x71_c, x72_c, x73_c, x74, x75, x77_c, x78_c, x79_c, x80_c, x81_c, x83, x84, x87_c, x88, x89_c, x90, x91_c, x92, x95, x96, x99);
and (w218, x8, x9_c, x14_c, x15_c, x21_c, x25_c, x31_c, x36_c, x39_c, x42_c, x46, x60, x61, x62, x67, x69_c, x73_c, x74_c, x75_c, x76, x77, x79_c, x83, x84, x85_c, x86_c, x88, x89_c, x90_c, x93_c, x95, x96, x97);
and (w219, x0, x7, x8, x12, x14, x28, x33_c, x34, x40_c, x41, x55, x58_c, x61_c, x62, x68_c, x72, x77, x80_c, x82, x84_c, x87, x92_c, x97_c);
and (w220, x0, x1_c, x2, x3, x4_c, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x13_c, x14, x15_c, x17, x18_c, x19_c, x20, x21_c, x22, x23, x24, x25, x26, x27, x28, x29_c, x30_c, x31, x32, x33, x34_c, x35, x36, x37_c, x39, x40_c, x41, x42_c, x43, x44, x45_c, x46_c, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57_c, x58, x59, x60, x61, x62, x63_c, x64, x65, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x72, x73, x74_c, x75, x76_c, x77, x78, x79, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87_c, x88_c, x89_c, x90, x91_c, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98_c, x99);
and (w221, x1_c, x3, x7_c, x8, x10, x11, x13_c, x16, x17, x21_c, x24, x26_c, x35, x45_c, x48_c, x49, x50, x52_c, x53, x56, x60_c, x62_c, x63_c, x64, x66_c, x75, x78_c, x85, x86_c, x93_c);
and (w222, x0, x4, x6_c, x7_c, x9_c, x12_c, x14_c, x16, x19_c, x22, x24_c, x25, x26_c, x27, x31, x35, x37_c, x38, x41_c, x42, x43_c, x44, x45_c, x46, x47, x49_c, x53, x55, x56_c, x61, x64_c, x65, x70_c, x71_c, x72, x74, x76_c, x77, x79_c, x82, x84, x87, x89_c, x90_c, x93_c, x94, x95_c, x96_c, x97_c);
and (w223, x0_c, x1, x3_c, x4_c, x5_c, x6_c, x7, x8, x9_c, x10_c, x11_c, x12_c, x14, x15_c, x16_c, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25, x26_c, x27_c, x28, x29, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50, x51, x52_c, x54_c, x55_c, x56_c, x57_c, x58_c, x59_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x70, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w224, x11_c, x13, x15_c, x18_c, x22_c, x26_c, x27_c, x30_c, x36, x37_c, x39, x42_c, x45, x50, x51_c, x54_c, x56, x60, x63_c, x66_c, x71_c, x72, x81, x85_c, x90_c, x97_c, x98_c);
and (w225, x8, x12, x18, x24_c, x27, x35_c, x39_c, x47_c, x51, x58, x62, x79, x80_c, x83);
and (w226, x2, x5_c, x6, x9_c, x12_c, x16_c, x24, x28, x31, x33, x36_c, x39, x40, x41, x42_c, x45_c, x49, x50, x55_c, x58_c, x59, x62, x64, x66, x70, x71, x73, x80_c, x83, x88_c, x92_c, x95);
assign w227 = x34;
and (w228, x3, x9_c, x14, x34_c, x37, x38_c, x47_c, x60, x67_c, x71, x75_c, x79_c, x81, x82_c, x91, x99_c);
and (w229, x0, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x33, x34, x35, x37, x38_c, x39, x41, x42, x43, x45, x46, x47, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68, x69, x70_c, x71, x72_c, x73_c, x74, x75, x77, x78_c, x79, x80, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x95, x96, x97, x98_c, x99_c);
and (w230, x4_c, x6_c, x12_c, x14, x20_c, x23, x31, x32, x33, x38, x39_c, x40, x42_c, x43_c, x44, x48, x53, x56, x58_c, x59, x60, x61, x63_c, x64_c, x66, x70, x72, x74, x75, x77, x78, x80_c, x82, x84_c, x87, x88, x94);
and (w231, x5_c, x11_c, x12, x13, x15, x16_c, x18, x20_c, x21, x23, x29_c, x31_c, x37, x51, x56, x57_c, x61_c, x70, x71_c, x76, x77, x82, x89_c, x90, x92, x94);
and (w232, x1, x3, x5_c, x49, x50_c, x64_c, x66_c, x70_c, x73, x79, x89, x92_c, x96);
and (w233, x0, x1_c, x2, x3, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x13_c, x14_c, x15_c, x16_c, x18_c, x19_c, x20_c, x21_c, x22_c, x24_c, x25, x26, x27, x28, x29_c, x30, x31_c, x32, x34_c, x36, x37, x38, x39_c, x40, x41, x44, x46_c, x47_c, x48_c, x49, x50_c, x52_c, x53, x54, x55_c, x56, x57, x59_c, x60, x61_c, x62, x63_c, x64, x65, x69, x70, x71, x74_c, x75_c, x76, x77_c, x78_c, x79_c, x81_c, x83, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92, x93, x94_c, x96_c, x97_c, x98_c, x99_c);
and (w234, x0, x3, x10, x13, x14, x15, x16_c, x22, x35_c, x38_c, x41, x46_c, x48_c, x52, x54, x58_c, x59, x64_c, x66_c, x74, x82_c, x84, x86_c, x91_c, x92_c, x93_c, x96_c, x97, x98);
and (w235, x0_c, x1_c, x2, x4, x6, x10, x11, x12_c, x13, x14, x15, x16, x17, x19, x20, x21_c, x22_c, x23, x24, x26_c, x27_c, x30_c, x31_c, x32, x34_c, x35, x37_c, x43_c, x47_c, x48_c, x49, x50_c, x51_c, x52_c, x53, x54, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x64, x65, x66, x69_c, x71, x72, x75, x77_c, x79, x81_c, x82, x83_c, x84_c, x85, x86, x88_c, x90, x91_c, x92_c, x93_c, x95_c, x96_c, x97, x98_c, x99);
and (w236, x1, x2_c, x3_c, x8, x10_c, x11_c, x16_c, x17_c, x18_c, x19_c, x20, x21_c, x22, x23, x25, x27, x28, x29, x30_c, x31_c, x32_c, x33_c, x35, x36_c, x37_c, x42_c, x43_c, x45_c, x46, x50_c, x54_c, x55, x60_c, x62, x63_c, x64, x66_c, x68, x69_c, x72, x73, x75, x78_c, x84, x85_c, x89_c, x90, x94, x96_c, x99);
and (w237, x0_c, x1_c, x2, x3_c, x4, x5, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14_c, x15, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30_c, x31_c, x32, x33, x34_c, x35, x37_c, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47_c, x48_c, x49_c, x50, x51, x52, x53_c, x55_c, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64, x65_c, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92_c, x93, x94, x95, x96, x97_c, x98_c, x99);
and (w238, x5, x7, x15_c, x23_c, x29_c, x38_c, x39, x40, x42, x44_c, x52, x53, x59_c, x65_c, x66, x74, x77_c, x81, x82, x87_c, x97);
and (w239, x0, x1, x2, x3, x5_c, x8_c, x9_c, x11, x12_c, x13, x14_c, x16, x18_c, x19_c, x20, x21_c, x22, x23, x24, x25_c, x26_c, x27, x28, x29, x30, x31_c, x32_c, x36_c, x37_c, x39_c, x41, x42_c, x43_c, x45, x47, x48, x49, x50, x51_c, x52_c, x54_c, x55, x58, x60_c, x62, x64, x65_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75, x76_c, x77_c, x79, x80_c, x81, x83_c, x84_c, x85, x86, x88, x89_c, x91_c, x92_c, x93_c, x94, x95, x96_c, x97_c);
and (w240, x40_c, x56, x92_c);
and (w241, x0, x1, x2, x3_c, x4, x5, x6, x7_c, x9_c, x10_c, x11, x12, x14, x17_c, x18_c, x19_c, x20_c, x21_c, x22, x23_c, x24, x25_c, x28_c, x29, x31_c, x35, x36, x37_c, x38_c, x39, x42, x43, x44, x46_c, x47, x48_c, x49_c, x50_c, x51, x52_c, x53_c, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x70_c, x72_c, x74, x75, x77, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x85_c, x86, x88_c, x89, x90, x92_c, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w242, x0_c, x1_c, x2, x3, x4, x5, x6_c, x7_c, x8, x9, x10_c, x12, x13, x14, x15, x16_c, x17_c, x18_c, x19, x20, x21, x22, x23, x24, x26_c, x27_c, x29, x30_c, x31_c, x32_c, x33, x34_c, x35, x36_c, x37, x38_c, x39_c, x40, x41, x42, x43, x44, x45, x46, x47, x48_c, x50, x51_c, x52_c, x53, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61, x62, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73_c, x74, x75, x76, x77, x78, x79_c, x80, x81, x82_c, x84_c, x85_c, x86_c, x87, x88_c, x89, x90, x91_c, x92_c, x93, x94, x95, x96_c, x98_c, x99_c);
and (w243, x0_c, x1, x3_c, x4, x5, x6_c, x7, x8_c, x9_c, x10, x12, x13, x14_c, x16_c, x17, x18_c, x19_c, x20_c, x21, x24, x26, x27_c, x28, x29_c, x32, x35, x36, x37, x45_c, x46, x49_c, x50_c, x52_c, x53, x55, x60, x65_c, x66_c, x67, x68_c, x69, x70_c, x72, x73_c, x75, x76, x78_c, x79_c, x81, x82_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92, x93, x94_c, x97_c, x98, x99);
and (w244, x0_c, x1, x2, x3, x4, x5_c, x6, x7, x8, x9, x10_c, x11, x12, x13_c, x15, x16, x17, x18, x19, x20, x21_c, x22, x25_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x33_c, x34_c, x35_c, x36, x37, x39_c, x40, x41_c, x42_c, x43_c, x44, x45_c, x46, x47, x48_c, x49, x51, x53_c, x54, x55_c, x57_c, x58, x59_c, x60_c, x61, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69_c, x70_c, x71, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x80, x81_c, x82, x84_c, x85_c, x86, x87, x88_c, x89_c, x90, x91, x92, x93_c, x95, x97, x98, x99_c);
and (w245, x1_c, x3, x4_c, x6, x7, x8_c, x10, x11_c, x12_c, x13, x15, x16, x18_c, x20_c, x21, x22, x23_c, x25, x26_c, x28, x34_c, x38, x40_c, x42_c, x43_c, x45_c, x46, x49_c, x53_c, x54, x56_c, x60_c, x61, x62, x63, x66, x67_c, x68, x69, x70_c, x72, x73, x75, x76, x78, x79_c, x82, x85, x86_c, x87, x91, x93, x94, x96, x99_c);
and (w246, x1_c, x2_c, x4, x5_c, x9_c, x10, x11_c, x13, x15_c, x16_c, x21, x23, x24, x25_c, x26, x28_c, x31, x34, x37_c, x42, x43, x46, x47, x48_c, x49, x50, x53_c, x54, x55, x56, x57, x59_c, x61_c, x64, x65, x70, x73_c, x75, x77_c, x78_c, x80, x81_c, x83, x85, x86, x90, x91, x94, x96);
and (w247, x11_c, x62, x69_c, x75, x92, x99);
and (w248, x0_c, x2_c, x3, x4_c, x5_c, x6, x7, x11_c, x13_c, x19_c, x20_c, x21_c, x22, x24, x27_c, x28_c, x29_c, x30, x32_c, x33, x34, x35_c, x36, x37_c, x38, x39, x40, x41_c, x42, x44_c, x46_c, x52_c, x54_c, x55, x57, x60, x62_c, x63, x65, x68_c, x69, x70_c, x71_c, x72_c, x73, x75, x78, x79, x80_c, x81_c, x83, x84, x86_c, x88_c, x89_c, x91, x92_c, x93_c, x95, x96, x97);
and (w249, x7_c, x12_c, x13, x25, x27, x31_c, x48_c, x49_c, x58, x59, x61_c, x62, x72_c, x73_c, x84_c, x87, x89_c, x90_c, x91_c);
and (w250, x7_c, x11, x19, x20, x21_c, x23, x28_c, x31_c, x35_c, x37, x39, x41_c, x42, x45_c, x47_c, x52, x53, x56_c, x68, x84_c, x90, x91, x92);
and (w251, x7, x9_c, x11_c, x40_c, x49, x54_c, x59, x66, x72, x74, x84_c, x86, x90, x92_c, x99_c);
and (w252, x0, x2_c, x3_c, x4_c, x5, x6_c, x7, x8, x9, x10, x11_c, x13, x14_c, x15, x16, x17, x19_c, x20, x21_c, x22, x23_c, x24, x25, x26_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35_c, x36, x37_c, x38, x39, x40_c, x43_c, x44, x45_c, x46_c, x47_c, x48_c, x49_c, x50, x51_c, x52, x53, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62_c, x63, x64, x65_c, x67, x68, x69_c, x70, x71, x73, x74_c, x75, x77_c, x78, x79_c, x80_c, x81_c, x82, x83, x84_c, x85_c, x87, x88, x89_c, x90_c, x91, x92, x93_c, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w253, x7_c, x12_c, x17_c, x19, x36_c, x41, x59, x64, x84, x91, x98_c, x99_c);
and (w254, x2, x6_c, x43_c);
and (w255, x4, x7, x8, x13_c, x15_c, x19_c, x20, x25_c, x27_c, x30, x35_c, x42, x43_c, x45, x46, x52, x56, x60, x61_c, x62_c, x70, x74_c, x75_c, x83, x87_c, x92_c, x94_c);
and (w256, x0_c, x1, x3_c, x5, x6_c, x8, x9, x10, x17_c, x18, x20_c, x21_c, x22, x24_c, x30, x31, x32, x33, x34_c, x37_c, x38_c, x42, x46, x47_c, x50, x53_c, x54_c, x55, x58, x59, x60, x61, x62, x63, x65, x66_c, x67, x69, x70, x71_c, x72, x73_c, x74, x75_c, x85, x87, x90, x91_c, x98_c, x99_c);
and (w257, x1, x3_c, x5, x9_c, x10_c, x13, x15_c, x17, x18, x19, x21_c, x22, x24_c, x25_c, x26, x27_c, x29_c, x30_c, x31_c, x32_c, x33, x39, x41_c, x42, x43_c, x44_c, x46, x47_c, x49, x50, x51_c, x53, x54, x55, x57, x58_c, x60, x61_c, x62_c, x65, x66, x67, x68_c, x69, x70_c, x71_c, x73_c, x75_c, x76, x77_c, x80, x81, x82_c, x86_c, x87_c, x88_c, x90_c, x91_c, x93_c, x95_c, x97_c, x98_c, x99);
and (w258, x2, x11_c, x31, x35, x42_c, x81, x97_c, x99_c);
and (w259, x5, x6_c, x13, x14_c, x18_c, x22, x29, x31_c, x34_c, x40_c, x47_c, x53_c, x59, x63, x70_c, x72_c, x73, x77, x78_c, x90_c, x96_c);
and (w260, x0, x2, x3_c, x4_c, x5_c, x8, x9_c, x10, x11_c, x12, x14_c, x15, x16, x17, x18_c, x19, x20_c, x21, x22_c, x23, x24, x25_c, x26_c, x27, x28_c, x29, x30, x33_c, x34, x37, x38_c, x41_c, x43, x44, x45, x46, x47, x48, x51, x52_c, x53, x54_c, x56, x57, x60_c, x61_c, x62, x63_c, x64_c, x65_c, x70_c, x71_c, x73_c, x76, x77, x82_c, x83_c, x84, x85_c, x86, x87, x92_c, x94, x95_c, x96_c, x97, x99_c);
and (w261, x0, x1, x2_c, x3, x4, x6, x7, x8_c, x9_c, x11_c, x12, x13, x14, x15_c, x17, x18, x19_c, x20, x21, x22_c, x23, x24, x25, x26, x27, x28, x29_c, x30, x31_c, x33_c, x34, x36_c, x37_c, x39, x40, x41, x42, x43, x44_c, x45_c, x46, x47, x48_c, x49, x50, x51_c, x52_c, x53_c, x54, x55_c, x56, x57, x58, x59_c, x60_c, x61_c, x62, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x80, x81_c, x82_c, x83_c, x84_c, x86_c, x87, x88_c, x89, x90_c, x92, x93_c, x94_c, x96, x97_c, x98, x99);
and (w262, x0, x1, x2_c, x4_c, x5, x6_c, x7, x8, x9, x11_c, x12, x13_c, x14_c, x15, x16_c, x17, x19, x20, x21_c, x22_c, x23, x25, x26, x27_c, x28, x29_c, x30, x31, x33, x34, x35, x37_c, x38, x40, x41_c, x42, x45_c, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62_c, x64_c, x65_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75_c, x76, x77, x81, x82_c, x83, x84, x85_c, x86, x88_c, x90_c, x91_c, x93, x94, x95_c, x96, x97_c, x98_c);
and (w263, x0_c, x1, x2_c, x3_c, x4_c, x5_c, x6, x7_c, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16, x17_c, x18, x19_c, x20, x21, x22_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x35, x36_c, x37, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46_c, x47, x48, x49_c, x50_c, x51, x52_c, x53, x54_c, x55, x56_c, x57, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65_c, x66_c, x67, x68, x69_c, x70_c, x71_c, x72, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80, x81_c, x82, x83_c, x84_c, x85, x86_c, x87_c, x88, x89, x91, x92_c, x93_c, x94_c, x95_c, x96_c, x98_c, x99_c);
and (w264, x1, x3_c, x7, x8_c, x9, x10_c, x12_c, x13_c, x14, x19_c, x21_c, x22_c, x24, x25, x27, x28_c, x30, x31_c, x36_c, x37_c, x38_c, x41, x42, x44, x47, x52_c, x53, x54_c, x55_c, x56, x59, x60, x65, x66_c, x73_c, x75_c, x78_c, x79_c, x81_c, x82_c, x83_c, x85, x86_c, x89_c, x90_c, x91, x99_c);
and (w265, x0, x1_c, x2, x3_c, x7, x8_c, x9_c, x10, x11, x12_c, x13, x14_c, x15_c, x17_c, x19_c, x20, x22, x23_c, x24_c, x25, x26, x27, x29_c, x30, x31_c, x32, x34, x35, x39, x40, x41, x42, x43, x44, x46_c, x47_c, x48, x49_c, x51, x52, x53_c, x54, x55_c, x56, x57_c, x58, x59_c, x60, x61_c, x62_c, x63, x64_c, x67_c, x68, x69, x70, x71, x72_c, x74_c, x75_c, x77_c, x78_c, x79, x80, x82, x83, x84_c, x85, x87, x88_c, x89, x91, x92, x94, x95_c, x96_c, x99_c);
and (w266, x0_c, x1_c, x3, x4_c, x9, x11, x13_c, x20, x23, x24_c, x26_c, x29_c, x30_c, x34_c, x38, x45_c, x46_c, x47_c, x48_c, x49, x51, x52, x56_c, x57, x59_c, x62, x64_c, x69_c, x70_c, x73, x74, x77, x80, x84_c, x89_c, x90, x97, x98_c);
and (w267, x3_c, x4_c, x5_c, x6_c, x7_c, x9_c, x11, x13, x15, x22_c, x23, x24_c, x25_c, x28, x31_c, x32, x34_c, x36_c, x40_c, x42_c, x43_c, x46_c, x49, x53_c, x54_c, x55, x58_c, x59_c, x72_c, x75_c, x76_c, x79_c, x80, x82_c, x84_c, x94, x99_c);
and (w268, x8, x12, x18_c, x20_c, x30_c, x31, x32, x33, x34_c, x37, x41_c, x43_c, x44, x46_c, x47_c, x49_c, x52, x53, x54_c, x55_c, x57, x63_c, x64, x65, x66, x67_c, x70, x73, x76_c, x77_c, x78, x82_c, x85_c, x86_c, x87, x93_c, x97_c);
and (w269, x1_c, x5, x9, x11_c, x12, x21, x24, x36, x37, x39_c, x41_c, x42_c, x43_c, x47, x48_c, x53_c, x55, x57, x58_c, x62_c, x67_c, x68_c, x70, x72_c, x74, x76, x77, x84, x85_c, x89, x93_c, x97_c, x98);
and (w270, x1_c, x2_c, x4_c, x5, x7_c, x8_c, x9_c, x10_c, x14, x15_c, x16, x17_c, x18_c, x20_c, x23, x25, x26_c, x28_c, x30, x31_c, x32, x37, x38, x44, x45_c, x47, x48, x52_c, x53, x54, x55, x57, x58, x59, x65, x66_c, x67_c, x68_c, x69_c, x71_c, x72, x73, x77, x79, x80, x81_c, x84, x85_c, x86, x87_c, x88, x90_c, x91_c, x92_c, x93, x96, x98, x99_c);
and (w271, x3, x5_c, x6, x7, x8_c, x13, x15_c, x16_c, x18_c, x19, x21, x22_c, x26, x28, x31, x33_c, x34, x38, x39_c, x42_c, x47_c, x48_c, x49_c, x50_c, x51, x53, x54, x56_c, x57, x58_c, x59_c, x62, x63, x66_c, x69_c, x70_c, x73, x74_c, x75, x76_c, x81, x83_c, x84, x87, x89_c, x90_c, x93_c, x94_c, x96, x99_c);
and (w272, x3_c, x5_c, x6, x7_c, x8_c, x10, x11_c, x12, x13_c, x14_c, x15, x16_c, x17, x18_c, x19_c, x22_c, x23, x24, x25_c, x27_c, x28, x29_c, x31, x33, x34, x35, x36_c, x38_c, x39, x40, x41_c, x42_c, x43_c, x44, x45_c, x46, x47_c, x49, x50_c, x51, x53, x54_c, x55, x57, x58_c, x59_c, x61_c, x62, x63, x64_c, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x71, x72, x74, x75_c, x76, x78, x79, x80, x81_c, x82_c, x84, x85, x86_c, x87, x88, x89_c, x90_c, x92_c, x93_c, x96, x98, x99);
and (w273, x2, x3, x8, x11, x12_c, x18, x22_c, x24, x40, x47_c, x50_c, x55, x60, x65_c, x70_c, x78, x81_c, x85_c, x86_c, x97_c);
and (w274, x0_c, x2, x3, x5, x6, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15_c, x16, x17_c, x18_c, x19_c, x20, x21, x22, x23, x25, x28_c, x29, x30, x31, x32, x33, x34_c, x35_c, x36_c, x37, x38, x39, x40, x41_c, x42_c, x43_c, x44, x46_c, x47_c, x48, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57_c, x58, x59, x60, x61, x62, x63_c, x64, x65, x66, x67_c, x68_c, x69_c, x71, x72_c, x73_c, x74_c, x75, x76_c, x78_c, x79_c, x80, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91_c, x93_c, x94_c, x96, x97_c, x98, x99);
and (w275, x0_c, x2_c, x3_c, x4_c, x6, x7, x8, x9_c, x10_c, x11, x12_c, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x24, x25, x26_c, x27, x28, x29, x30_c, x31_c, x32, x33, x34, x35, x36_c, x38, x40_c, x41, x42, x43, x44, x45_c, x46_c, x47, x48_c, x49, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57, x58_c, x59, x60, x61, x62, x63_c, x64_c, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x74, x75, x76_c, x77_c, x79, x80, x81_c, x82_c, x83, x84, x86_c, x88_c, x89, x90, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w276, x0, x1, x3, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x13_c, x14, x15, x16_c, x17, x18_c, x20, x22_c, x23, x25_c, x29, x33_c, x35, x36_c, x38, x39_c, x41_c, x42, x43, x44, x45_c, x46, x47_c, x48_c, x54, x55, x58_c, x59, x60_c, x63, x68, x69_c, x70, x73_c, x74_c, x75_c, x76_c, x77, x79_c, x81, x82, x84_c, x92_c, x96_c, x98, x99_c);
and (w277, x1, x2_c, x3, x4, x5, x6, x7_c, x8_c, x9_c, x11, x13_c, x14, x15, x16_c, x17, x19_c, x20, x21, x22_c, x23, x24, x26, x27_c, x29_c, x30_c, x31_c, x32_c, x33_c, x38_c, x40_c, x41_c, x43_c, x45, x47, x48_c, x49_c, x50, x52_c, x53_c, x54, x55_c, x60, x61_c, x63, x64, x67, x69_c, x70, x71, x73, x74, x75_c, x77, x78_c, x80_c, x81_c, x82, x83_c, x84_c, x85_c, x88_c, x89_c, x90, x91_c, x92_c, x93, x99);
and (w278, x1, x3, x4_c, x8_c, x9, x10_c, x13, x15_c, x16_c, x18_c, x19_c, x20_c, x23_c, x24_c, x25_c, x26_c, x27_c, x29_c, x31, x33_c, x36_c, x37_c, x38_c, x40, x43_c, x45_c, x46, x47, x48, x49_c, x51, x52_c, x53, x54_c, x55_c, x56, x61, x62_c, x63_c, x65, x66_c, x67, x68_c, x71_c, x72_c, x73_c, x75, x76_c, x77_c, x78, x79_c, x80_c, x82, x83, x84, x85, x86_c, x87, x88, x90_c, x91, x92_c, x93, x94, x95, x96, x97, x98);
and (w279, x1, x2, x3_c, x4, x5_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13, x14_c, x15, x16_c, x17_c, x18_c, x19, x20, x22_c, x23, x24, x25, x26_c, x27, x28, x29_c, x30_c, x31_c, x33_c, x34, x36, x37, x38_c, x39, x40_c, x41_c, x42, x43_c, x44, x45_c, x46, x47_c, x48, x49_c, x51, x52, x53_c, x54_c, x56, x57_c, x58_c, x59, x60_c, x61_c, x62_c, x63, x64_c, x65, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x73_c, x75_c, x76, x77, x78_c, x79_c, x80, x81, x82_c, x83_c, x84, x85_c, x86_c, x87, x88, x89_c, x90_c, x91, x92_c, x93, x94, x96, x97, x98_c);
and (w280, x0, x1_c, x2, x3, x4, x6, x7_c, x8_c, x9, x10_c, x12, x13, x14, x16_c, x17, x18_c, x19_c, x20_c, x21, x22_c, x23, x24_c, x26, x27, x28_c, x29_c, x30, x31_c, x32, x33_c, x36_c, x37, x38_c, x41, x42, x43_c, x44, x46, x47, x48_c, x49_c, x50, x51, x52, x53_c, x54_c, x55_c, x58_c, x59_c, x60_c, x62_c, x64, x65_c, x67_c, x68, x70_c, x71, x72, x73, x74_c, x75, x76_c, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x88, x89, x90, x91, x93_c, x95_c, x96, x97, x99);
and (w281, x1_c, x3_c, x4_c, x5_c, x6, x9_c, x10, x11_c, x13, x17, x20, x22_c, x23, x25_c, x26_c, x28, x29_c, x30_c, x31, x35, x37_c, x40, x42_c, x43_c, x49, x51, x52_c, x53, x54, x57_c, x58_c, x59_c, x61, x62_c, x64, x66, x67_c, x69, x70, x71, x72_c, x73, x75, x80_c, x81_c, x85, x86_c, x88_c, x89, x93_c, x95_c, x96, x98_c, x99_c);
and (w282, x1_c, x3_c, x4_c, x5_c, x6, x7, x8_c, x9, x10, x11_c, x13, x14, x16, x18, x19_c, x20, x21, x22_c, x23, x24, x25, x26_c, x27_c, x28, x30, x31_c, x32, x33_c, x35, x36_c, x37_c, x38_c, x40, x41_c, x42_c, x43, x44_c, x45_c, x46, x47_c, x48_c, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56_c, x57_c, x58_c, x59_c, x60, x62, x63_c, x64, x65, x66, x67, x69, x70, x71, x72, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x81, x82, x83_c, x84, x87_c, x88, x89_c, x91, x92_c, x94_c, x95, x96, x97, x98_c, x99_c);
and (w283, x0_c, x1_c, x2, x4, x5, x8, x9, x10_c, x11, x13, x14_c, x15_c, x17_c, x18, x20_c, x21, x22, x23_c, x26_c, x27, x28, x29_c, x30_c, x33, x35, x36, x37_c, x38, x39, x40_c, x41_c, x44, x45_c, x46, x49_c, x50_c, x52, x53_c, x54, x56_c, x57, x58, x60, x61_c, x62_c, x65_c, x66, x69, x72_c, x73, x74, x75_c, x79, x81_c, x85, x87, x88_c, x91_c, x93, x95_c, x96, x97_c, x98, x99_c);
and (w284, x0, x1, x2, x3, x4, x5, x6, x7_c, x8, x9, x10_c, x12, x13, x15, x16, x17, x18, x19_c, x20_c, x21_c, x22, x23_c, x25_c, x26, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x41_c, x42_c, x43, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51_c, x52_c, x53_c, x54, x55, x56_c, x57, x58_c, x59, x60, x61_c, x62_c, x63, x64_c, x65, x66, x67_c, x68_c, x69, x70, x71, x72_c, x73, x74_c, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x82, x83_c, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97, x98_c, x99_c);
and (w285, x0, x1_c, x11, x12, x14_c, x15_c, x17, x19, x20_c, x21_c, x22_c, x24, x28_c, x29_c, x30_c, x31_c, x32, x34, x35, x36, x37, x39, x40_c, x41_c, x42, x44, x45, x46_c, x47_c, x48_c, x51, x52, x53_c, x56_c, x57, x58, x59_c, x62_c, x63_c, x65, x66_c, x67_c, x69_c, x70, x73, x75, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83, x84, x85_c, x87_c, x90, x91_c, x92_c, x93_c, x94, x96);
and (w286, x0, x2_c, x3_c, x4_c, x5_c, x6, x7, x9, x12_c, x14, x16, x17, x18, x19, x20_c, x21, x26_c, x28_c, x29, x35, x38, x41, x42_c, x43_c, x46_c, x47, x48, x51, x52, x53, x54_c, x55_c, x56, x58, x59_c, x60_c, x63_c, x64_c, x65, x66_c, x68_c, x71, x72, x73_c, x74_c, x77, x78_c, x79_c, x81_c, x83_c, x86, x90_c, x91, x93, x95, x97, x98);
and (w287, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7_c, x8, x9_c, x10, x11, x12, x13_c, x14_c, x15, x16_c, x17_c, x18_c, x19, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x34, x35, x36, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55_c, x56_c, x57_c, x58, x59_c, x60, x61_c, x62, x63_c, x65_c, x66_c, x67, x69_c, x70_c, x71_c, x72, x73_c, x75_c, x76_c, x77, x78, x79, x80, x82_c, x83_c, x84_c, x85, x86_c, x87_c, x88, x89_c, x90, x91, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w288, x0, x1_c, x5, x6_c, x7, x8, x12, x13_c, x18, x25_c, x33_c, x36, x37_c, x39, x41, x46_c, x48, x49_c, x51_c, x55_c, x62, x68_c, x70, x71_c, x72_c, x74_c, x75, x76, x77, x79_c, x81_c, x86_c, x88_c, x89, x90, x91, x92, x94, x95_c, x98_c);
and (w289, x0, x1, x2_c, x3, x5, x7_c, x8, x9, x10_c, x12_c, x14_c, x15_c, x16_c, x17, x18, x20_c, x21_c, x22, x23_c, x25, x26, x27_c, x28_c, x29, x30, x32, x34_c, x35_c, x36, x37_c, x38_c, x39, x40, x42, x43, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50_c, x51, x52_c, x53_c, x54_c, x56, x57_c, x58_c, x59, x60_c, x62_c, x63, x64, x65, x67, x68, x69_c, x70, x71, x72_c, x73_c, x75, x76, x77_c, x78_c, x79_c, x81_c, x82, x83, x84, x86, x87, x88_c, x89, x90_c, x91_c, x92_c, x93, x95, x96, x97_c, x98);
and (w290, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x8, x10_c, x11_c, x12, x13_c, x14_c, x16, x17_c, x18, x19_c, x20, x21_c, x22_c, x23, x24, x25_c, x27, x28_c, x31, x32, x33, x34, x35_c, x36_c, x37, x38, x39_c, x40, x41_c, x43, x45_c, x46_c, x48_c, x49_c, x50_c, x51, x53_c, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62_c, x65_c, x66_c, x67_c, x70, x71, x72_c, x74, x76, x77_c, x78_c, x80_c, x81_c, x82, x83_c, x84_c, x85_c, x86, x87_c, x88_c, x89, x90, x92_c, x93_c, x97_c, x98_c, x99_c);
and (w291, x0_c, x1_c, x2_c, x3_c, x4_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x15, x16_c, x17, x18_c, x19_c, x20_c, x21, x22, x23, x24, x25, x26, x28_c, x30, x31, x32_c, x33, x34, x35, x36, x37, x38, x39_c, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48_c, x49_c, x50, x51, x52, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x63, x64, x65, x66, x67_c, x70, x71, x73_c, x74, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x83, x85, x86, x87, x88_c, x89_c, x90_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99_c);
and (w292, x2_c, x5, x23, x24, x39, x60, x66, x68_c, x70, x84_c);
and (w293, x5_c, x7_c, x10, x13, x14_c, x16, x19, x20_c, x21_c, x22, x25, x27, x33, x42_c, x45, x47_c, x48, x49_c, x54_c, x58_c, x60, x66_c, x71, x72_c, x73_c, x77_c, x82_c, x85_c, x86, x87, x91, x92, x94, x95);
and (w294, x0, x1_c, x2, x3_c, x4, x5, x6_c, x7_c, x9, x10, x12_c, x13_c, x14, x15_c, x16, x19_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x40_c, x41_c, x42_c, x43, x45_c, x47, x48_c, x51_c, x52, x53_c, x54_c, x56, x58_c, x59, x60_c, x61, x62, x63, x66, x67_c, x69, x74, x75, x76_c, x77_c, x78, x79, x80_c, x81, x83_c, x84, x88, x89, x92, x94_c, x95_c, x96_c, x97_c, x99_c);
and (w295, x0_c, x2_c, x8, x9_c, x10_c, x11, x13, x14_c, x15, x16, x17_c, x18_c, x19, x21, x25, x27_c, x28_c, x29_c, x30, x31_c, x34_c, x35, x36_c, x37_c, x38, x39, x41, x42_c, x43_c, x44, x45_c, x46_c, x49, x50, x51_c, x52, x53, x54_c, x55_c, x56_c, x58, x60_c, x63, x64_c, x65, x66, x67, x69, x71_c, x72, x73_c, x74, x75, x77_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x86_c, x89, x90_c, x92, x93_c, x98);
and (w296, x5, x8_c, x10_c, x11, x14, x21, x22_c, x28, x32_c, x33, x47, x49_c, x51, x57, x63, x67_c, x74_c, x77, x80_c, x84, x88, x94);
and (w297, x0, x4_c, x12_c, x22_c, x27_c, x30, x32_c, x39, x43_c, x48, x54, x69_c, x78_c, x92, x96);
and (w298, x32_c, x51, x60);
and (w299, x0_c, x1, x2_c, x3_c, x4, x6, x7, x8, x9_c, x10, x11, x12, x14_c, x16_c, x17, x19, x21_c, x22_c, x24, x25_c, x26_c, x27, x28, x29_c, x30, x31_c, x33_c, x34, x35, x36, x37_c, x38, x39_c, x40, x42, x43, x44, x45_c, x46, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x57, x58, x59_c, x60_c, x62, x63, x64, x66_c, x67, x68_c, x70_c, x71, x72_c, x73, x74_c, x75_c, x77, x78, x82_c, x83, x84_c, x85_c, x86, x87, x88, x89, x91_c, x92, x94_c, x96_c, x97, x98_c, x99);
and (w300, x2, x8_c, x10, x14, x16, x22_c, x23, x24, x27, x29_c, x31, x32, x33, x36, x38_c, x40, x42_c, x45_c, x46_c, x50, x59, x63, x68_c, x76, x85_c, x87_c, x89, x91, x95, x97_c, x98_c);
and (w301, x0_c, x2, x3, x4, x5, x6, x7, x10_c, x11, x12, x13, x14_c, x15_c, x16_c, x17_c, x18, x19_c, x21, x23_c, x24, x25_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36_c, x37, x38_c, x39, x40, x42, x43_c, x44, x45, x46, x48_c, x49, x50, x51, x52, x53, x54, x55_c, x57, x58_c, x59_c, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70, x71, x72, x74_c, x76_c, x77, x78, x79, x80_c, x81_c, x83, x84, x85_c, x86, x88, x89_c, x90, x91, x92, x93, x94, x95_c, x96, x97_c, x98, x99);
and (w302, x1, x2_c, x4_c, x6, x7_c, x8_c, x11, x14_c, x17, x18_c, x20, x21_c, x22, x23, x24, x25_c, x26, x27_c, x29_c, x30_c, x32, x35_c, x37, x38_c, x42_c, x44_c, x45_c, x47_c, x48_c, x50, x52, x53_c, x54, x56, x57_c, x58_c, x62_c, x63, x65, x66_c, x67, x68_c, x69, x70_c, x72_c, x74, x77_c, x78_c, x79, x80_c, x82_c, x85, x86_c, x87_c, x88, x89_c, x90, x91, x92_c, x95_c, x96);
and (w303, x1, x27_c, x35, x36_c, x45, x48, x50, x58, x86_c, x87_c, x92_c);
and (w304, x2_c, x4_c, x10, x16, x20, x21, x22_c, x29, x31_c, x32, x40, x45, x47, x50, x53_c, x55, x56, x57_c, x59_c, x61_c, x63, x65_c, x66_c, x70_c, x73, x74, x75, x78_c, x80_c, x87_c, x88, x98, x99);
and (w305, x0, x1, x2, x5, x6_c, x7, x12, x14, x15, x16_c, x17_c, x19, x22_c, x23, x25, x26, x27, x29_c, x30, x31_c, x32, x33, x34_c, x36_c, x39, x40_c, x41_c, x44, x45_c, x47_c, x48_c, x49, x51_c, x52_c, x54, x56, x57, x58_c, x59_c, x60_c, x61_c, x62_c, x66, x67_c, x68_c, x70, x71_c, x72, x73_c, x74_c, x76_c, x78, x79, x80, x81_c, x82_c, x83, x85_c, x86, x87_c, x88, x90, x91_c, x92, x93_c, x94_c, x97_c, x98, x99);
and (w306, x0, x3_c, x4, x6_c, x7, x8, x9_c, x11_c, x12, x13_c, x15, x17, x18_c, x19_c, x22_c, x23, x24_c, x25_c, x26, x28, x30, x31_c, x33_c, x35, x38, x40, x42_c, x43_c, x45, x46_c, x47, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x55, x57_c, x58, x59, x60, x61_c, x62, x64_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x72, x73_c, x74, x75, x76_c, x77, x80, x81_c, x83_c, x84, x88, x90_c, x92_c, x95_c, x98_c);
and (w307, x2_c, x3_c, x5, x7, x8_c, x9, x10_c, x11_c, x12_c, x13, x14_c, x16_c, x21_c, x23, x24_c, x25, x26_c, x28_c, x29, x30, x31_c, x32, x33, x34, x35_c, x37_c, x38, x39_c, x40_c, x41, x42, x43, x44_c, x45, x46_c, x47_c, x48_c, x51_c, x53_c, x54, x56, x57_c, x58_c, x59, x60, x61, x62_c, x63_c, x66_c, x68_c, x69, x70, x71_c, x72_c, x73, x74, x75, x76, x77_c, x79_c, x80, x81, x83_c, x84, x86_c, x87_c, x89, x90_c, x91, x92_c, x93_c, x95, x97, x98_c, x99_c);
and (w308, x0, x2, x3_c, x4, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11, x13_c, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22_c, x23, x24, x25_c, x26_c, x27, x28_c, x30, x31_c, x32_c, x33, x34_c, x35, x36, x37, x38, x39, x40, x41_c, x42_c, x43, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50, x51, x52_c, x53_c, x54_c, x55, x58_c, x59, x61, x62_c, x63_c, x64, x65, x66, x67, x68, x69_c, x70, x71, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78, x79, x80_c, x81, x82_c, x83, x86, x87_c, x88_c, x89, x90, x91_c, x92, x93_c, x94, x95, x96_c, x97_c, x98, x99);
and (w309, x0_c, x1, x2, x4_c, x5_c, x6_c, x8_c, x9_c, x10, x11, x12, x13_c, x14, x15, x16_c, x17_c, x18, x19, x20_c, x21, x22, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35_c, x37_c, x38, x39_c, x40, x41_c, x43, x44_c, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52, x53, x55, x56_c, x57, x58_c, x59, x60_c, x61, x62_c, x63, x64_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71_c, x72, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83, x84, x85, x86, x87, x88_c, x89_c, x90_c, x91_c, x92, x93_c, x94_c, x95_c, x96_c, x97, x98, x99_c);
and (w310, x3, x6, x8_c, x10, x12_c, x14_c, x16, x19_c, x25, x34, x35_c, x38_c, x39_c, x40_c, x41, x42, x45_c, x46_c, x47_c, x48, x51, x53_c, x56_c, x59, x60_c, x63_c, x65_c, x70, x73, x75, x76, x77, x78, x79, x81, x83_c, x86_c, x89_c, x95_c, x97_c);
and (w311, x0, x2, x11_c, x19_c, x20_c, x30_c, x34_c, x37_c, x40_c, x54, x57_c, x62_c, x78, x79, x80_c, x95, x99_c);
and (w312, x26_c, x28_c, x40_c, x44, x57_c, x62, x71_c);
and (w313, x0_c, x1, x5, x6, x7, x8_c, x10, x11, x13, x18_c, x22_c, x23_c, x24, x27, x33, x34, x35_c, x40_c, x41, x42, x43, x46, x49_c, x52, x54, x56, x57_c, x59, x60, x63_c, x64_c, x66, x68, x69, x71, x72_c, x73_c, x74_c, x75_c, x77, x79, x81, x83, x84, x86_c, x87_c, x93_c, x94, x95_c, x96, x97_c, x98_c, x99_c);
and (w314, x0_c, x1, x2_c, x5, x10, x11_c, x13, x16_c, x17, x19, x22, x24, x25_c, x26_c, x32, x33_c, x38, x40_c, x41, x42_c, x46_c, x47, x49, x51, x52_c, x53, x56_c, x58_c, x59, x62, x63, x64_c, x66_c, x69, x70, x72, x73_c, x76, x77, x84_c, x86_c, x90_c, x94_c, x95, x96_c, x97_c, x99);
and (w315, x0_c, x6, x8_c, x10_c, x11, x12_c, x13_c, x14, x15_c, x16_c, x17, x18_c, x22_c, x23, x28_c, x31, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39_c, x41, x43_c, x49, x51, x52_c, x53, x54, x55_c, x57_c, x60, x61_c, x62, x63_c, x66, x67, x70_c, x72, x74, x75, x77_c, x79_c, x80, x82_c, x84, x85, x86, x87_c, x89_c, x96_c, x97);
and (w316, x39_c, x88_c);
and (w317, x0_c, x2_c, x6_c, x7, x8_c, x10_c, x11_c, x12_c, x14, x15, x17_c, x18, x19, x21, x22_c, x23, x25_c, x26, x27, x29_c, x30, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x42_c, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50_c, x51, x55, x56_c, x57_c, x58, x59_c, x60_c, x61, x62, x63_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x74_c, x75, x77_c, x78_c, x79_c, x81_c, x83_c, x84_c, x85, x87, x89, x91, x92, x93_c, x95_c, x96, x97, x98_c, x99);
and (w318, x23, x39, x55_c, x64, x65, x70, x74);
and (w319, x0, x4_c, x5_c, x6_c, x7_c, x8_c, x11, x16_c, x18_c, x19, x22, x23, x26, x27, x28, x29, x33, x34, x36, x37_c, x40_c, x41_c, x42_c, x44_c, x46, x47, x49_c, x50, x51, x52_c, x53_c, x54, x56, x57, x60, x61, x63_c, x64, x65_c, x67, x68, x69_c, x70, x72, x75, x76, x77, x79_c, x80_c, x81_c, x83_c, x85, x86_c, x88_c, x91_c, x92, x93, x96, x97, x98_c);
and (w320, x20_c, x25, x31, x35, x51_c, x68);
and (w321, x12_c, x14);
and (w322, x3_c, x5_c, x6_c, x7, x8_c, x9, x14_c, x15, x17_c, x18, x19_c, x21_c, x22, x23, x25, x26_c, x27_c, x28, x30_c, x31_c, x32, x33, x35_c, x36, x38_c, x39_c, x41_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48, x49_c, x50, x52, x53_c, x54, x55, x56, x57_c, x58_c, x59, x60_c, x62, x63_c, x64_c, x65_c, x67_c, x68, x69, x70, x71, x72_c, x73_c, x74_c, x76, x77, x78, x79_c, x80, x81_c, x82, x83_c, x84, x86, x87_c, x88_c, x89_c, x90_c, x92, x94, x95, x96, x97, x98);
and (w323, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x8_c, x9, x11, x12, x13_c, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x23_c, x24_c, x25_c, x27, x28, x29_c, x30, x31, x32, x33_c, x34, x35, x37, x38_c, x40, x41, x42_c, x43, x45, x47, x48_c, x49, x50_c, x51, x52, x53, x54, x55_c, x56_c, x58, x59_c, x61, x62, x63, x64, x65, x67_c, x68, x69_c, x70_c, x71, x72, x73_c, x75, x76_c, x77, x78, x79_c, x80, x81, x82_c, x83, x84_c, x85, x86, x87, x89, x91, x93, x94, x95_c, x96, x97, x98_c);
and (w324, x11_c, x43, x53_c, x78, x90_c);
and (w325, x0, x2_c, x3, x5_c, x6, x9, x14_c, x15, x16, x18_c, x19, x20_c, x24, x26, x27, x28_c, x31, x39, x43, x47, x48, x50, x51, x65, x68_c, x69_c, x71_c, x72_c, x73, x74_c, x79, x80_c, x81, x86_c, x87, x96, x97, x99);
and (w326, x0, x1, x2_c, x8, x9_c, x10, x17, x21, x26_c, x27_c, x29_c, x34_c, x40, x41_c, x42_c, x45_c, x48, x49, x50, x54_c, x56, x59, x62, x65_c, x66, x68_c, x75_c, x78_c, x80_c, x82, x85_c, x89_c, x92, x93, x94, x95, x96, x97, x98, x99_c);
and (w327, x0, x2, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x20_c, x21_c, x22, x23_c, x25_c, x26_c, x29_c, x30_c, x31, x33_c, x37_c, x40_c, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x51, x53, x56_c, x57, x58, x60_c, x61, x62_c, x65, x66, x67_c, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x79_c, x83, x85, x86_c, x87, x90_c, x92_c, x93_c, x94, x95, x96, x99_c);
and (w328, x7, x9, x15, x17, x21_c, x24_c, x29, x34, x37_c, x42_c, x46, x50_c, x51, x55_c, x63, x64, x66, x67, x68, x69, x72_c, x73, x79_c, x83_c, x89, x92_c, x93, x97_c, x98, x99);
and (w329, x1, x7, x8, x10_c, x16, x20, x22_c, x29_c, x36, x39, x45, x47, x51_c, x52_c, x55, x57, x60, x61, x66_c, x72, x74, x75_c, x91_c, x98);
and (w330, x0, x2, x4, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x22_c, x24_c, x25_c, x26, x29, x30_c, x33, x34, x35_c, x36_c, x37_c, x40_c, x41_c, x46_c, x48, x51, x52_c, x53_c, x54_c, x55_c, x57_c, x59, x60_c, x64_c, x65, x68_c, x70_c, x71_c, x72_c, x73_c, x74, x77, x78, x79_c, x81, x82_c, x83_c, x84, x85, x87_c, x89, x91, x92_c, x97, x98, x99_c);
and (w331, x2, x9_c, x14, x21, x29_c, x36_c, x50, x70_c, x93, x96_c);
and (w332, x0, x1, x2, x3_c, x4_c, x5_c, x6, x7, x8_c, x9, x10, x11, x12, x13, x14, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27, x28, x29, x30, x31_c, x32, x33, x34, x35, x36, x37_c, x38_c, x39, x40, x41_c, x42, x43, x44, x45_c, x46, x47, x48, x49_c, x50, x51, x52_c, x53, x54_c, x55_c, x56, x57, x58_c, x59, x60_c, x61, x62, x63_c, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73_c, x74, x75, x76, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90_c, x91, x92_c, x93, x94_c, x95, x96_c, x97_c, x98, x99);
and (w333, x1_c, x17, x19_c, x30_c, x42_c, x43, x44_c, x55, x56, x59, x64_c, x66_c, x73, x82_c, x86_c, x90_c);
and (w334, x5, x7, x10_c, x11, x12, x15_c, x20_c, x22_c, x27_c, x29_c, x31_c, x35_c, x39, x50_c, x60, x68_c, x71_c, x79, x84_c, x88, x90, x93);
and (w335, x0_c, x3, x5, x7_c, x8, x9_c, x10, x11, x12, x13_c, x14_c, x15_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x25, x26, x28, x29_c, x30, x31_c, x32, x33, x34_c, x35_c, x36, x37_c, x39, x40_c, x42, x43, x44, x45_c, x46, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61, x62, x63, x64_c, x65, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x73, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83_c, x84, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92, x93_c, x94_c, x95_c, x96_c, x98_c, x99);
and (w336, x33, x34_c, x36_c, x40, x41_c, x63, x66_c, x67, x71_c, x94_c, x97_c);
and (w337, x2, x3_c, x4_c, x15, x24, x34, x36_c, x39_c, x41_c, x42_c, x47, x52, x54, x56_c, x57, x68, x69_c, x70, x81, x82, x86_c, x92, x97_c, x99);
and (w338, x0, x1_c, x3, x4, x5, x6, x8_c, x9, x10_c, x11, x12, x13_c, x15_c, x16, x17_c, x18, x19_c, x24, x25, x26, x27_c, x28, x29_c, x30_c, x32_c, x33, x34_c, x35_c, x36, x37, x38, x39_c, x40, x41_c, x42_c, x45_c, x46_c, x47, x49_c, x50, x51_c, x52, x53_c, x54, x55_c, x56_c, x58_c, x59, x60, x61, x62, x63, x64_c, x65, x67, x68, x69, x70, x71_c, x72_c, x73, x74_c, x76_c, x77_c, x78_c, x79_c, x80, x82, x83_c, x84_c, x85, x87, x88, x89_c, x90, x92, x93, x94_c, x96_c, x97, x98, x99);
and (w339, x0, x1_c, x2_c, x3_c, x5_c, x6, x7, x8_c, x9, x10_c, x11, x12, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24, x25, x26, x27, x28, x29_c, x30, x31, x32_c, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x54, x55_c, x56_c, x58_c, x59_c, x60, x61, x63_c, x64, x65, x66, x67, x68, x69_c, x70, x71_c, x72, x73, x74, x75, x76, x77, x78_c, x79, x80, x81_c, x82_c, x83_c, x84, x85_c, x86, x87, x88, x89, x90_c, x91_c, x92, x93_c, x94, x95, x96, x97_c, x98_c, x99_c);
and (w340, x0, x1, x3, x4, x5_c, x6, x7_c, x8_c, x9_c, x10, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23, x24_c, x25, x26, x27_c, x28_c, x29_c, x30_c, x31_c, x32, x33, x34_c, x35, x36, x37_c, x38, x39_c, x40_c, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x50, x51_c, x52, x53, x54, x55_c, x56, x57_c, x58, x59, x60, x61, x62, x63, x64, x65_c, x66_c, x67, x68, x69, x70, x71, x72, x73, x74_c, x75, x76, x77_c, x78, x79, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92, x93, x94, x95, x96, x97_c, x98, x99_c);
and (w341, x0_c, x3_c, x10, x15, x16_c, x19_c, x20_c, x22_c, x23, x27, x29, x30, x33, x34, x35, x42, x43_c, x53_c, x57_c, x60_c, x62_c, x63, x64_c, x69, x71_c, x72_c, x75, x77, x79, x80, x85, x86_c, x93, x96_c);
and (w342, x1_c, x3_c, x7_c, x8, x9_c, x10_c, x11_c, x12, x16_c, x17, x18_c, x23_c, x25_c, x26_c, x27, x30_c, x31, x32_c, x33_c, x40, x42, x44_c, x45_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52, x55, x56_c, x57, x58_c, x61_c, x62_c, x65_c, x66_c, x69_c, x70, x72, x73_c, x75_c, x77, x79_c, x80_c, x81, x86, x88, x90, x91, x92_c, x96_c, x97_c, x99_c);
and (w343, x0_c, x1_c, x2_c, x3, x4, x6, x7, x8, x9_c, x10, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17, x18, x19, x20_c, x21, x22_c, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x38_c, x39_c, x40_c, x42, x44, x45, x46_c, x49, x51_c, x52_c, x53, x54, x55, x57, x58_c, x59, x60_c, x61, x62, x63, x64, x66, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x75_c, x76, x77_c, x78_c, x80, x81_c, x82_c, x83_c, x84_c, x85, x86, x87_c, x88, x89, x90, x91, x93, x94_c, x95, x96_c, x97, x98_c, x99_c);
and (w344, x0_c, x4, x17, x57, x75_c, x83, x90_c);
and (w345, x1, x4, x6, x8_c, x9_c, x10, x11, x13_c, x14, x15, x16, x18, x19_c, x20_c, x21_c, x22, x24, x25_c, x26, x27, x30, x31_c, x32_c, x36_c, x39_c, x40_c, x41_c, x42_c, x43, x46_c, x48, x49_c, x50_c, x52_c, x54, x55, x57_c, x58, x59, x63, x64_c, x67_c, x70, x71_c, x72_c, x74, x77, x79_c, x81, x82_c, x83, x84_c, x87_c, x88, x89_c, x91, x93_c, x94, x95, x98, x99_c);
and (w346, x0, x5_c, x6, x10_c, x11_c, x15, x17, x18, x19_c, x20_c, x21_c, x22, x27_c, x29_c, x30_c, x32, x33_c, x34, x36_c, x37, x42, x45_c, x46_c, x48_c, x50_c, x54, x59, x60_c, x61_c, x62, x69, x70, x73, x74_c, x78_c, x80, x81, x83_c, x85_c, x86, x90, x91_c, x92, x95_c, x97_c, x99);
and (w347, x0, x3, x4, x8_c, x9, x10_c, x12, x16, x17, x20_c, x23_c, x24, x25, x26, x27_c, x28, x29_c, x30_c, x33, x35_c, x36, x38_c, x40_c, x41_c, x42_c, x44, x45_c, x46_c, x50_c, x51_c, x52, x53, x54, x55_c, x56, x58_c, x59_c, x63_c, x65, x66, x67_c, x68_c, x70_c, x73_c, x76, x78, x79, x80_c, x82_c, x84, x85, x89, x90, x92_c, x93_c, x94_c, x96_c, x98);
and (w348, x0_c, x2_c, x4_c, x7, x8, x14_c, x15_c, x17, x21_c, x23_c, x28_c, x29, x31, x36_c, x40_c, x41, x46, x48, x52, x53, x57_c, x59_c, x62, x63_c, x64_c, x67, x68_c, x74_c, x77_c, x78_c, x79_c, x81, x82_c, x83_c, x84_c, x88_c, x96_c);
and (w349, x20_c, x28_c, x32, x40, x41, x43, x44, x49_c, x52, x55_c, x60_c, x65_c, x71, x72, x73_c, x75, x84, x85_c, x89_c, x92, x93, x98, x99_c);
and (w350, x0, x41_c, x58_c, x60_c, x63, x83_c, x85);
and (w351, x0, x1_c, x2_c, x3, x4_c, x5_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23, x24, x25_c, x26, x27, x28, x29, x30, x31, x32_c, x33_c, x34_c, x35, x36_c, x37, x38_c, x39_c, x40, x41_c, x42, x43_c, x44_c, x45, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57_c, x58, x59, x60, x61_c, x62, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78, x79, x80, x81, x82_c, x83_c, x84, x85_c, x86, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x97, x98, x99);
and (w352, x9, x13, x17, x19, x28_c, x37, x42, x47_c, x54, x64_c, x85, x86, x89_c, x91_c, x93_c, x96);
and (w353, x1, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11, x12, x13_c, x15_c, x16_c, x17, x18_c, x19, x20, x21, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31, x32_c, x33_c, x34_c, x35_c, x36, x37_c, x38_c, x39, x40, x41, x42, x44_c, x45, x46, x47, x48_c, x49, x50, x51_c, x52, x53, x54, x55, x56, x57_c, x58, x59_c, x65_c, x67_c, x68_c, x69, x70_c, x71, x72, x73_c, x74, x76_c, x77, x78_c, x79, x80_c, x81_c, x82, x83_c, x85_c, x86_c, x87, x88_c, x89_c, x90, x91_c, x92, x93_c, x95, x97, x98);
and (w354, x1, x5, x7_c, x17, x18, x19, x20_c, x22, x23, x24_c, x31_c, x32, x35_c, x38, x40_c, x41, x43, x47_c, x49_c, x53_c, x54_c, x57, x58_c, x59, x76, x79_c, x80_c, x81_c, x85, x89_c, x90_c, x91, x99);
and (w355, x0, x1, x2, x4_c, x5_c, x6_c, x7, x11_c, x12_c, x13, x15, x16_c, x17_c, x18, x19, x20, x23_c, x24, x26, x28_c, x29_c, x30_c, x31, x32, x34_c, x35_c, x36_c, x37, x38, x39_c, x41, x42_c, x43, x46_c, x47_c, x48, x50_c, x51_c, x52, x53_c, x54, x56, x57_c, x58_c, x60, x61_c, x63, x64_c, x65, x66, x67, x68_c, x71_c, x72, x74, x75_c, x76_c, x77_c, x79_c, x83, x84_c, x86_c, x87, x88, x89, x91_c, x92_c, x94, x95, x96_c, x98, x99_c);
and (w356, x8_c, x11, x19, x43_c, x44_c, x50_c, x69, x81_c);
and (w357, x0_c, x1, x2_c, x3, x4, x7, x8_c, x9, x10, x11, x12, x13_c, x14_c, x15, x16_c, x17_c, x18, x19_c, x20_c, x21, x22_c, x23, x24_c, x25_c, x26_c, x28, x29, x30_c, x31_c, x32, x33, x34, x35, x36, x37, x38, x39_c, x40, x41_c, x43, x44_c, x45_c, x47_c, x48_c, x49, x50, x51_c, x52_c, x53, x54_c, x55, x56, x57_c, x59, x60_c, x61, x63, x65, x66_c, x67, x69, x70, x71, x72_c, x73, x74, x76_c, x77, x78, x80, x81, x83_c, x84, x85_c, x86, x87, x88, x89_c, x90, x91, x92, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w358, x0, x1, x2_c, x4_c, x5, x6_c, x8, x9, x10_c, x11, x12_c, x14, x15, x17_c, x18_c, x20_c, x21_c, x22, x23, x24_c, x25, x27, x28, x30, x32, x33, x34_c, x35, x37_c, x38, x40, x41, x42, x43_c, x44_c, x45, x46_c, x47_c, x48, x49, x50, x51, x52, x53_c, x54, x55_c, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64, x66_c, x67_c, x69, x70, x71, x74_c, x75_c, x76, x79, x80, x81_c, x83_c, x86, x87_c, x89_c, x90_c, x92, x93, x94, x95_c, x97, x98_c, x99_c);
and (w359, x0, x1, x2, x5, x6_c, x7_c, x9_c, x11, x13_c, x14_c, x17, x18_c, x19_c, x20, x21, x22, x27_c, x29_c, x32, x33, x36, x38, x40, x41, x42_c, x43_c, x45_c, x46, x49_c, x50_c, x51_c, x52_c, x55_c, x57, x58_c, x60_c, x61_c, x63_c, x64, x65_c, x67, x69_c, x72_c, x74, x75_c, x77, x78, x79_c, x80, x81, x82, x83_c, x86_c, x90, x91_c, x92, x94_c, x96_c, x97, x99_c);
and (w360, x0_c, x1_c, x2, x3, x5, x6_c, x7, x9_c, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x20_c, x21, x22, x24, x27_c, x29_c, x33, x34_c, x35_c, x36_c, x37, x40_c, x41, x42, x44_c, x45, x46, x49_c, x50, x51_c, x52, x54, x56, x57_c, x58_c, x59, x60, x62_c, x64_c, x65, x69, x70, x71_c, x72_c, x73, x75_c, x77, x78_c, x79, x81, x82, x83, x86_c, x87_c, x89, x91, x92_c, x96_c, x97);
and (w361, x6_c, x9, x29, x66_c, x69_c, x81_c, x82_c, x94_c);
and (w362, x7, x8, x15, x18, x20, x21_c, x26_c, x27, x28, x34, x42, x45_c, x47, x50, x51_c, x52_c, x56_c, x58_c, x69, x71, x76_c, x79, x82, x83_c, x87_c, x92, x94, x96_c, x97_c);
and (w363, x12, x13, x14, x16_c, x19, x22, x27, x30_c, x44, x56, x71_c, x98_c);
and (w364, x30_c, x64);
and (w365, x0, x1_c, x3, x4_c, x6_c, x8_c, x12_c, x14, x20_c, x23, x24_c, x26_c, x29_c, x31_c, x32_c, x34, x36, x38, x40, x41_c, x43, x47, x52_c, x55_c, x58, x64_c, x66, x70, x74_c, x78_c, x79_c, x81, x84_c, x86_c, x92, x94, x98_c, x99);
and (w366, x0_c, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8_c, x9, x10_c, x13_c, x14_c, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x29_c, x30_c, x31, x34, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x45, x47, x49_c, x50_c, x51, x52_c, x53, x54, x55, x56, x57, x58_c, x61_c, x64_c, x65_c, x66, x67_c, x69, x70_c, x73_c, x74_c, x78, x79, x81, x83_c, x84, x85, x86_c, x87, x89, x93_c, x95_c, x96_c, x97_c, x99_c);
and (w367, x1_c, x3_c, x4, x10_c, x12_c, x13_c, x15_c, x36, x38_c, x39, x42_c, x43_c, x48, x52_c, x57, x58_c, x59, x60_c, x63, x65_c, x68_c, x76, x82, x86_c, x99_c);
and (w368, x3_c, x4, x5, x8, x9_c, x10_c, x12_c, x17, x18_c, x19, x20_c, x21, x22, x23_c, x24, x26, x28, x29_c, x30, x31, x35, x37, x42_c, x45_c, x47_c, x48, x50_c, x51_c, x53, x55, x56, x57_c, x58_c, x59, x61, x62, x63, x65_c, x66_c, x67_c, x69, x73_c, x74_c, x75_c, x76, x79, x82_c, x85_c, x86_c, x89, x93);
and (w369, x0_c, x4_c, x7, x8_c, x12, x13_c, x14_c, x18_c, x19_c, x21, x37_c, x38, x46_c, x47, x48, x49_c, x52_c, x53, x55_c, x57, x58_c, x61, x63, x66_c, x67, x68_c, x72, x75_c, x83, x84, x86, x87_c, x89, x91, x97_c);
and (w370, x3_c, x8_c, x18, x27_c, x45, x49_c, x50, x51, x53_c, x56, x68_c, x83_c, x84, x89, x92_c);
and (w371, x0_c, x1_c, x3, x5, x6_c, x7_c, x8_c, x9, x10, x11_c, x12_c, x13_c, x14_c, x19_c, x21, x22, x23, x26_c, x27_c, x28, x29, x30, x31, x33_c, x34, x35, x36_c, x38_c, x39_c, x40, x41_c, x44_c, x45_c, x48, x49, x51, x52, x54_c, x55_c, x56_c, x57_c, x58_c, x60_c, x62, x63_c, x64_c, x66, x67_c, x69, x70, x72, x73_c, x74_c, x76, x77_c, x79, x82, x89_c, x90_c, x91, x92, x94_c, x96_c, x98);
and (w372, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16, x17_c, x18_c, x19_c, x20, x21, x22_c, x23_c, x24_c, x25, x26_c, x27_c, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x35, x36_c, x38, x39_c, x41, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x54, x55_c, x56_c, x57_c, x58_c, x59, x60, x61, x62, x63_c, x64_c, x65, x66_c, x68, x69, x70_c, x71, x72, x73_c, x74_c, x77, x79_c, x80, x81_c, x82, x83_c, x86_c, x87_c, x88_c, x89, x90, x91_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w373, x0_c, x2_c, x5, x7, x8_c, x11, x13, x14_c, x16, x18_c, x19, x20, x21_c, x22, x23, x24_c, x25, x26_c, x27, x29_c, x35_c, x36_c, x40_c, x42, x46_c, x48_c, x49, x58, x59, x60, x61, x62, x63, x64, x65_c, x66_c, x67, x68_c, x69_c, x70_c, x75_c, x76_c, x77_c, x79_c, x82_c, x83, x84_c, x87, x88, x90_c, x91, x92, x93, x94_c, x98);
and (w374, x6, x13_c, x21_c, x24_c, x34, x46_c, x51, x57_c, x60, x61_c, x62, x65_c, x68, x74, x92_c, x94_c);
and (w375, x0, x1, x2_c, x3, x4_c, x5_c, x6, x7_c, x8, x9_c, x10_c, x11_c, x12, x14_c, x15, x16_c, x17_c, x18_c, x19, x20_c, x21, x22, x24, x25, x26_c, x27_c, x28, x30, x31, x33_c, x34_c, x35_c, x37_c, x38, x39_c, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x49_c, x50_c, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61, x62, x66_c, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80_c, x81, x82_c, x83, x84, x85_c, x86_c, x87, x88_c, x89, x90_c, x92, x93_c, x94, x95, x97, x98_c, x99);
and (w376, x0_c, x1, x2, x3, x4_c, x5, x6, x7, x8_c, x9, x11, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22_c, x23_c, x24_c, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34, x36_c, x37, x38, x39_c, x41, x42_c, x43_c, x44, x45, x46, x47, x48, x50_c, x51, x52_c, x53_c, x54_c, x55, x57, x58_c, x59, x62_c, x63_c, x64, x65_c, x66, x67, x68_c, x69_c, x70, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x90_c, x91, x92, x93_c, x94, x95_c, x96, x98_c, x99);
and (w377, x1_c, x3_c, x7, x8, x9, x10, x11_c, x12_c, x13_c, x14, x18, x20_c, x21, x25_c, x26, x27_c, x28_c, x29, x30, x33, x38, x43, x44, x45_c, x48, x50_c, x51, x52_c, x53_c, x55, x58, x61_c, x62_c, x63_c, x64_c, x66_c, x67, x68, x70_c, x71, x72, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x82_c, x84, x85_c, x87, x89_c, x92_c, x93_c, x94_c, x95, x97, x99);
and (w378, x1_c, x2, x4_c, x6_c, x7, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14, x17, x21, x22_c, x24_c, x26_c, x28, x29_c, x32_c, x33, x34_c, x35, x37_c, x38, x39, x42, x43_c, x44, x45, x49, x50, x51_c, x53_c, x54_c, x55_c, x58, x59_c, x60_c, x61_c, x62, x63_c, x64, x65, x66, x67_c, x68_c, x70, x71, x72_c, x73, x74_c, x75_c, x76, x78, x80, x81_c, x82, x83_c, x85, x86, x88_c, x89_c, x95, x96_c, x98_c, x99);
and (w379, x0_c, x1, x2, x3, x4_c, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12, x13, x14, x15, x16, x17_c, x18, x19_c, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30_c, x31, x32, x33, x34, x35_c, x36_c, x37, x38, x39, x40_c, x41, x42, x43, x44_c, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51, x52_c, x53_c, x54_c, x55_c, x56_c, x57, x58_c, x59_c, x60_c, x61, x62_c, x63, x64_c, x65, x66, x67_c, x68_c, x69_c, x70, x71_c, x72, x73, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81_c, x82_c, x83, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96_c, x97, x98, x99);
and (w380, x2_c, x8_c, x25_c, x27, x36_c, x45_c, x47, x62, x72, x73, x75_c, x91, x99_c);
and (w381, x16_c, x18_c, x19_c, x20, x22, x26, x32_c, x35, x40, x44_c, x46, x47, x53, x55, x58, x61_c, x64, x65, x68, x71_c, x72, x75, x78, x81_c, x83, x89_c, x90, x94_c, x95_c, x98);
and (w382, x0_c, x1, x3_c, x4, x6_c, x8, x9_c, x11_c, x13_c, x15_c, x17_c, x19_c, x21, x23, x24_c, x28_c, x29_c, x30_c, x31, x32_c, x33, x34, x36, x39, x41, x42_c, x47_c, x49_c, x50_c, x54, x56_c, x58, x59_c, x60, x61_c, x62_c, x63_c, x64, x65_c, x70, x73_c, x74, x75, x77, x80, x81, x83_c, x84_c, x87, x88, x89, x91, x92_c, x93, x95_c, x97_c, x98_c);
and (w383, x6, x13, x18, x20, x22_c, x31, x34_c, x38, x44_c, x46_c, x47_c, x54, x58, x61, x64, x68_c, x71_c, x74_c, x75_c, x76_c, x79, x80, x81, x99);
and (w384, x0, x1, x3_c, x4, x5, x7, x10_c, x13, x14, x15, x17, x18_c, x19, x22, x23_c, x24_c, x28_c, x30, x32_c, x33_c, x37_c, x38, x40, x41, x44_c, x46, x47_c, x53, x57_c, x59_c, x68_c, x71, x74_c, x75, x77_c, x78, x79, x82, x83_c, x89, x90_c, x93, x96_c, x97_c);
assign w385 = x23_c;
and (w386, x0, x1_c, x2_c, x3, x4, x5, x7, x9, x10_c, x12_c, x13, x15_c, x17, x18_c, x21_c, x23_c, x25, x26, x27_c, x28, x29_c, x31, x32, x33, x34_c, x35, x38, x39_c, x40, x43, x44_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54, x55, x56, x57, x59, x60, x61, x62, x63_c, x64, x66, x67_c, x69, x71, x72_c, x73_c, x75_c, x76, x77, x78, x79, x80, x81_c, x87_c, x89_c, x90_c, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w387, x0_c, x1, x2, x4_c, x5, x6, x7, x8, x9_c, x10, x12, x13_c, x14, x15, x17_c, x18, x19_c, x20, x21_c, x24, x25, x26, x27_c, x28, x30_c, x32, x33, x34, x35_c, x36, x39_c, x42, x43, x45_c, x46_c, x47_c, x48_c, x50_c, x51_c, x53_c, x54_c, x56_c, x57, x58, x59, x60, x61_c, x62_c, x65_c, x66_c, x68, x69, x70, x71_c, x73_c, x74, x75_c, x76_c, x77, x79, x80_c, x81, x82_c, x83, x84, x85, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x94_c, x95_c, x96_c, x97, x98, x99);
and (w388, x0, x1, x2_c, x3, x4, x5_c, x6, x7, x8, x9_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29, x30, x31_c, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x39_c, x40, x42_c, x43, x44, x45_c, x46, x47, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x56, x57, x58_c, x59_c, x60, x61_c, x62, x63, x64_c, x65_c, x66_c, x67, x68, x69_c, x70, x71_c, x72_c, x73, x74_c, x75, x77_c, x78, x79, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x89_c, x90, x91, x93_c, x94_c, x95_c, x96, x97, x98);
and (w389, x13_c, x14_c, x37_c, x39_c, x45_c, x53_c, x54, x55, x67_c, x78, x82, x83);
and (w390, x1, x4, x11_c, x12, x14_c, x16, x17_c, x20_c, x36, x41_c, x43_c, x44_c, x46_c, x48_c, x49_c, x52, x53_c, x54, x56_c, x59, x62, x71_c, x77_c, x79_c, x80, x83_c, x86_c, x89, x90_c, x91, x95, x96);
and (w391, x0_c, x2_c, x3_c, x4_c, x6, x7_c, x8, x9_c, x10_c, x11, x12, x13_c, x14, x16, x17, x19_c, x20, x21, x22, x23, x25_c, x27, x31_c, x33, x34, x36_c, x37, x39, x40, x42_c, x43, x44, x45_c, x46_c, x47_c, x48, x49, x50_c, x51_c, x52_c, x55, x56_c, x57, x64_c, x65_c, x66, x67_c, x68, x74, x76, x77_c, x78_c, x79, x80, x81, x84_c, x85, x88_c, x89_c, x93_c, x94_c, x96, x97, x99_c);
and (w392, x0_c, x3_c, x7, x9, x11, x17, x21_c, x24, x32_c, x36_c, x38, x43, x44, x45_c, x47_c, x53, x58_c, x61, x62, x65_c, x69, x73, x81_c, x84_c, x87_c, x91_c, x92);
and (w393, x0, x2_c, x4, x10, x12, x13_c, x16, x23_c, x24, x25_c, x32, x33_c, x35, x36_c, x41, x49_c, x50_c, x53_c, x56_c, x62, x63_c, x65_c, x67_c, x74_c, x75_c, x82, x84_c, x87, x88_c, x92, x93, x94_c, x97);
and (w394, x2, x4_c, x6_c, x7_c, x12_c, x13, x20, x23_c, x35, x36_c, x47, x50, x51, x70_c, x78_c, x90_c, x96);
and (w395, x13, x14, x23, x24_c, x29_c, x30_c, x42, x43_c, x45, x53_c, x55_c, x56, x64_c, x76_c, x80);
and (w396, x3_c, x12_c, x16_c, x20, x44_c, x52, x66, x69_c, x92_c);
and (w397, x0_c, x1_c, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15_c, x16, x17_c, x18, x20, x21, x23_c, x25, x26_c, x27, x29, x30, x32_c, x33_c, x35, x36, x37_c, x39, x41_c, x42, x43, x45_c, x47_c, x49, x50_c, x51_c, x55, x56, x57, x58_c, x62, x63_c, x64, x65, x66, x68_c, x69, x70, x71, x72_c, x73_c, x75, x77_c, x78_c, x79_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x91_c, x93, x95_c, x96_c, x98_c, x99_c);
and (w398, x0_c, x1_c, x2_c, x3, x4_c, x5, x6_c, x9, x10_c, x13_c, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x27, x28, x29, x30_c, x31_c, x33, x34, x35_c, x36, x37, x38_c, x39, x40_c, x41_c, x42_c, x44_c, x45, x46, x47, x48_c, x49_c, x53_c, x54, x55, x56, x57_c, x58, x59_c, x60, x61_c, x64_c, x67_c, x68_c, x69_c, x70_c, x72, x73, x74_c, x76, x77_c, x78, x79, x81, x82_c, x83_c, x84, x85, x86, x88_c, x89_c, x92_c, x93_c, x94, x95_c, x96_c, x99_c);
and (w399, x0, x1, x2, x3, x5, x9, x10, x12_c, x13_c, x14, x15, x17_c, x18_c, x21_c, x22_c, x24_c, x25, x26_c, x29, x30_c, x31_c, x32, x33, x36, x37_c, x38_c, x39, x41_c, x42_c, x43, x44_c, x45_c, x48_c, x49_c, x53, x54, x58, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69, x70, x71_c, x72, x74, x75_c, x76, x78_c, x79, x80, x81_c, x82, x83_c, x85, x87, x88_c, x89, x90_c, x91_c, x92_c, x93, x94_c, x95, x98_c);
and (w400, x1, x3, x5_c, x6_c, x8_c, x9, x10_c, x11_c, x12, x13, x16_c, x18_c, x19, x21_c, x22, x23, x25_c, x26_c, x27_c, x28_c, x30, x31, x34, x36_c, x37_c, x38_c, x39, x40_c, x41_c, x42, x43_c, x44, x47_c, x48, x50_c, x51, x55_c, x57, x58_c, x59_c, x60, x63, x64, x65_c, x66, x69, x70_c, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x80, x81_c, x82, x83_c, x84_c, x85, x88_c, x89, x90, x91_c, x92_c, x94, x95, x96, x97_c, x98);
and (w401, x0_c, x5, x23_c, x30_c, x31, x32, x38_c, x42_c, x46, x47, x50_c, x51, x54_c, x56_c, x61_c, x63_c, x65, x72_c, x81, x84, x85, x95);
and (w402, x0, x1_c, x2_c, x4, x6_c, x8_c, x13, x14_c, x17_c, x20, x23_c, x27, x28_c, x29, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x39_c, x46_c, x47_c, x48_c, x50, x51, x52, x53, x54, x55_c, x57, x59_c, x61_c, x62, x63_c, x64_c, x66, x68, x69, x70_c, x71, x73_c, x74, x75, x77_c, x78_c, x79, x80_c, x83, x84_c, x87, x92_c, x93, x94_c, x95, x99);
and (w403, x0_c, x1_c, x4_c, x5, x6_c, x8, x10_c, x12_c, x13_c, x15, x16_c, x18, x22_c, x23, x25, x26_c, x27_c, x32_c, x36_c, x37, x38, x39, x40_c, x41_c, x43_c, x44, x45, x46, x47, x48_c, x51, x53, x54_c, x55_c, x57_c, x58_c, x60_c, x63, x65_c, x69_c, x70, x71_c, x72, x76_c, x77_c, x78_c, x80, x81_c, x82, x83_c, x85, x87_c, x96_c, x97_c);
and (w404, x0, x1, x2, x3, x5, x6, x7, x8, x9_c, x10_c, x11, x13_c, x14_c, x15_c, x16_c, x17_c, x18_c, x19, x20_c, x23_c, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31, x33_c, x34_c, x35_c, x36_c, x37, x38, x39_c, x40_c, x42, x43_c, x44, x45, x46_c, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x57, x58_c, x59_c, x60_c, x61_c, x62_c, x64_c, x65_c, x67_c, x68_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77, x78, x79_c, x80_c, x81, x82_c, x84, x85_c, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94, x95, x96_c, x98, x99_c);
and (w405, x3, x21_c, x26_c, x29, x39, x40, x55, x79, x83, x96_c, x97);
and (w406, x0_c, x1, x2, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x11, x12, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21, x22, x23, x24_c, x25_c, x26, x27, x28_c, x29_c, x30, x31_c, x32_c, x33, x34_c, x35, x36_c, x37_c, x38_c, x39_c, x40, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50_c, x51_c, x52_c, x53_c, x54, x55, x56, x57, x58, x59, x60, x61_c, x62, x63, x64, x65, x66_c, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85_c, x86, x87, x88_c, x89, x90, x91, x92, x93, x94_c, x95_c, x96_c, x97, x98, x99_c);
and (w407, x0, x1, x4, x5_c, x6, x7, x8_c, x9_c, x10, x11_c, x12_c, x13, x15_c, x16, x17, x18, x19_c, x20, x21, x22_c, x23_c, x24_c, x25, x27_c, x29_c, x30_c, x31, x32, x33, x35_c, x36_c, x38, x40_c, x41, x42, x43, x45, x46_c, x47, x48, x49, x50_c, x51, x54, x55, x56_c, x57_c, x59_c, x60_c, x61, x62_c, x63, x64_c, x65, x66, x67, x69_c, x70, x72, x73_c, x75_c, x77, x78_c, x79, x81, x82, x83_c, x84, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93_c, x95, x97_c, x98);
and (w408, x0_c, x2_c, x14_c, x17, x18, x28, x30_c, x33, x36, x37_c, x40, x45_c, x49_c, x50, x60, x69_c, x71, x72, x75_c, x82, x85, x97);
and (w409, x6_c, x7, x8_c, x12_c, x13_c, x14_c, x26_c, x32, x35, x42, x48_c, x49, x55_c, x57_c, x58_c, x66_c, x69_c, x77_c, x79_c, x82, x97_c);
and (w410, x0_c, x1, x2_c, x3_c, x5_c, x7_c, x8_c, x11_c, x12, x14_c, x15, x16_c, x17_c, x20_c, x23_c, x24_c, x25, x26_c, x28_c, x29, x32, x34, x35, x36, x37_c, x38, x40_c, x42, x43, x44_c, x45, x47_c, x48_c, x49, x50_c, x51_c, x52, x56_c, x57_c, x58, x61, x62, x68_c, x69_c, x71, x74, x76, x77_c, x78_c, x79, x80_c, x81_c, x83, x84_c, x86, x87_c, x88, x89_c, x90, x92_c, x94, x95, x96_c, x97_c, x98_c, x99_c);
and (w411, x0, x1, x2_c, x3, x4, x5_c, x6, x7, x8_c, x11_c, x16_c, x17, x18, x19, x20_c, x21, x22_c, x24, x25, x28, x30_c, x31_c, x32_c, x33, x34, x35_c, x36_c, x40_c, x41, x42_c, x43, x44, x45, x46, x47, x48, x50, x51, x52_c, x54, x56_c, x60, x61_c, x63_c, x65_c, x66, x67_c, x68_c, x70, x72, x73, x76, x82, x83_c, x85_c, x86, x88, x89, x92_c, x93_c, x94, x95, x96, x97, x99);
and (w412, x0_c, x1, x2, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29, x31_c, x32, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45, x46, x47_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x64, x65_c, x69, x70_c, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x87_c, x89, x90_c, x91, x93, x94_c, x95, x96, x97);
and (w413, x0, x26_c, x30_c, x36_c, x37, x48, x74_c, x96);
and (w414, x5_c, x9, x27, x61_c, x76, x88_c);
and (w415, x5, x10, x16, x21_c, x34_c, x35, x41, x42_c, x45, x73_c, x76, x85, x89);
and (w416, x0_c, x2_c, x4, x6, x8_c, x11_c, x13_c, x16_c, x17_c, x18_c, x19, x21_c, x22_c, x23, x24_c, x28, x29, x32_c, x33_c, x34, x35, x36, x37, x38_c, x39, x40, x41_c, x43, x45, x46_c, x47, x48, x49, x50, x51_c, x53_c, x55_c, x56_c, x59_c, x60_c, x61, x62, x64, x65, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x73, x75, x76_c, x77, x78_c, x81, x82, x83_c, x84_c, x85, x87, x89, x90_c, x91, x92, x93, x94_c, x95_c, x96_c, x97, x98, x99);
and (w417, x2_c, x8_c, x9_c, x32, x33_c, x37_c, x39_c, x40, x54_c, x56_c, x57, x68_c, x70, x75, x79, x87, x89, x91_c, x94, x97);
and (w418, x2_c, x3, x4_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x14_c, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x39_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x50, x51_c, x52, x53_c, x54, x55, x56, x59, x60, x61_c, x62_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x76_c, x78, x79_c, x80, x81_c, x82, x83_c, x84_c, x85, x86, x89, x90, x91_c, x93_c, x94_c, x95_c, x96, x97_c, x98_c, x99_c);
and (w419, x0, x1_c, x3, x4, x5_c, x7, x10, x12, x14_c, x15_c, x16, x17, x18, x20_c, x22, x23, x24_c, x25, x28, x29, x30_c, x31_c, x32, x33_c, x34_c, x35_c, x37, x38, x39_c, x40, x42_c, x43_c, x44, x46, x47, x49, x50, x51, x52_c, x57_c, x58_c, x60_c, x61, x62_c, x63_c, x65_c, x67_c, x68, x69_c, x70, x71, x72, x73_c, x74, x75_c, x77_c, x78_c, x80, x81, x82_c, x84_c, x85, x86, x87_c, x88_c, x89_c, x90, x91_c, x93_c, x94, x96, x97, x98_c);
and (w420, x3_c, x8_c, x14, x23_c, x24, x29, x31, x36, x47_c, x53_c, x58, x69, x74, x78_c, x80_c, x86, x87_c, x88, x89, x90, x98_c);
and (w421, x0_c, x1, x2_c, x3_c, x4_c, x5_c, x6, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23, x24_c, x26_c, x27, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35_c, x36, x37, x39_c, x40, x41, x42_c, x43, x44_c, x45_c, x46_c, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x57, x58, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w422, x3_c, x5, x8, x15, x16_c, x19, x20_c, x21_c, x25_c, x26_c, x28, x31_c, x32, x33_c, x35_c, x36, x37, x44, x47_c, x48, x50, x56_c, x59_c, x64_c, x67, x68, x77_c, x80_c, x81, x86, x90, x91_c, x92, x94_c, x96, x98);
and (w423, x0_c, x2_c, x3_c, x7_c, x16, x38_c, x40_c, x42_c, x51, x72, x90, x93, x97);
and (w424, x33_c, x52, x99_c);
and (w425, x0_c, x1_c, x2_c, x5_c, x6_c, x7, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18, x19_c, x20, x21_c, x22_c, x23_c, x24_c, x25, x26, x27_c, x28_c, x29_c, x31_c, x33, x34_c, x35, x36_c, x37_c, x39, x41_c, x45_c, x46, x48, x49_c, x50_c, x52_c, x53_c, x54, x55_c, x56_c, x57, x59_c, x60_c, x63_c, x64, x66, x67, x70_c, x71_c, x72, x73, x74_c, x75, x76, x77, x78, x79, x81_c, x82_c, x83_c, x84_c, x86, x88, x90_c, x92_c, x93, x94, x96_c, x97_c, x98);
and (w426, x0, x1_c, x2_c, x3_c, x4, x5_c, x6, x7, x8_c, x9_c, x10, x11_c, x12_c, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24, x26_c, x27, x28_c, x29, x30, x31, x32_c, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54_c, x56_c, x57, x58_c, x59, x60_c, x61, x62, x63, x64, x65, x66_c, x67, x68_c, x69, x70, x71_c, x72_c, x73_c, x74_c, x75_c, x76, x77_c, x78, x79, x80, x81, x82, x83, x84_c, x85_c, x86, x87, x88, x89_c, x90_c, x91, x92_c, x93_c, x94_c, x95, x96_c, x97, x98, x99_c);
assign w427 = x29;
and (w428, x1, x12_c, x21, x51, x64, x74_c, x78_c, x96_c);
assign w429 = x23_c;
and (w430, x2, x3, x6, x7, x8, x9, x12_c, x14_c, x16, x17, x24_c, x25_c, x26_c, x29, x32, x34_c, x35_c, x39_c, x40_c, x41_c, x42_c, x48_c, x49_c, x50, x53, x55, x56_c, x62, x63_c, x64, x65, x69_c, x70, x71_c, x72, x74, x75_c, x76_c, x77, x80_c, x81_c, x83_c, x84, x85_c, x88, x91, x92, x94_c, x96, x97, x98);
and (w431, x0_c, x1_c, x2, x3, x4, x6, x7_c, x8, x9_c, x10, x11, x12_c, x13_c, x14_c, x15, x16, x17_c, x18, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x34, x35, x36, x37, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45_c, x46, x48_c, x49, x50_c, x51_c, x52_c, x53, x54, x56, x57_c, x58_c, x59, x60, x61_c, x62_c, x63_c, x65, x66, x68, x69, x70_c, x71, x72_c, x73, x75, x76, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85, x86, x87_c, x88, x89, x90, x91, x93_c, x94_c, x95, x96_c, x99_c);
and (w432, x2_c, x3_c, x4, x6, x7, x8, x10, x11, x14, x16, x17, x19, x21, x25, x27, x28, x30_c, x31, x32_c, x35_c, x36_c, x37_c, x39, x40, x42, x43_c, x44, x45, x46_c, x49, x50, x52_c, x54, x57, x58_c, x59, x60, x62, x65, x66, x68_c, x69_c, x72_c, x73_c, x82, x83, x84_c, x88_c, x89, x91_c, x92, x93, x97, x98);
and (w433, x2_c, x6_c, x8, x10_c, x11_c, x14_c, x17, x18_c, x22_c, x24, x25_c, x31, x33_c, x38_c, x41, x47, x49_c, x50_c, x52, x58, x60, x62_c, x65_c, x71_c, x74, x75_c, x77, x78_c, x81, x84, x89_c, x95_c, x96);
and (w434, x0, x2, x3_c, x4, x6_c, x7_c, x10, x11_c, x18, x19, x20_c, x21, x24, x25_c, x26_c, x27_c, x28, x30_c, x32_c, x33, x35_c, x37, x39, x40_c, x42_c, x43_c, x46_c, x47_c, x48, x49, x52, x54_c, x55, x56_c, x58_c, x59, x61_c, x62_c, x63, x67_c, x69_c, x70_c, x72, x73, x74_c, x75_c, x77, x78_c, x79, x80_c, x81, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x92_c, x94_c, x95_c, x96_c, x97_c);
and (w435, x0, x1_c, x2_c, x3, x5, x6_c, x7, x8_c, x9_c, x10_c, x11_c, x13_c, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x21, x23_c, x24, x25_c, x26, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34, x35, x36_c, x37_c, x38, x39, x40_c, x41, x42_c, x43, x44_c, x45_c, x46, x47_c, x48, x49, x50_c, x51, x52, x53, x54, x55, x56, x57, x58_c, x59, x60, x61, x62, x63, x64, x65_c, x67, x68, x69_c, x70_c, x72_c, x73_c, x75_c, x77, x78_c, x80_c, x81, x82, x83, x84, x85, x86, x87_c, x88_c, x90_c, x91, x92, x93, x94, x95_c, x97, x98, x99_c);
and (w436, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8, x10_c, x11_c, x12, x13, x14_c, x15_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x44, x45, x46, x47_c, x51, x52_c, x53, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70_c, x71, x72, x73, x74_c, x75_c, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94, x95, x96_c, x97, x98);
and (w437, x0, x1_c, x2, x3, x4, x6_c, x7_c, x8, x9, x10_c, x11_c, x12, x15_c, x18, x20, x21, x23, x27_c, x28_c, x30_c, x37, x41_c, x42_c, x44, x46_c, x49, x57, x60_c, x61_c, x64, x66, x71_c, x72, x73_c, x76_c, x77_c, x78, x82, x83_c, x95_c, x96, x97_c, x98, x99_c);
and (w438, x0_c, x1_c, x2_c, x3, x4_c, x5, x6_c, x7, x8, x9, x10_c, x11, x12, x13_c, x14, x15, x16, x17, x18, x19_c, x20_c, x21_c, x22, x23, x24, x25, x26, x27_c, x28, x29, x31, x32, x33, x34_c, x35_c, x36, x37_c, x38, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x46, x47_c, x49_c, x50_c, x51, x52, x53_c, x54, x55, x57, x58, x59_c, x60, x61_c, x62_c, x63, x64, x65_c, x66_c, x67, x68_c, x69, x70, x71, x72_c, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x90, x91, x92_c, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w439, x0_c, x2, x3_c, x4, x6_c, x7, x9, x10, x14_c, x15, x17, x18, x29_c, x31_c, x32, x33_c, x34, x35, x40_c, x43_c, x44, x46_c, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x56_c, x57, x58, x59_c, x60, x61_c, x62_c, x63, x64, x65_c, x66_c, x67, x68, x69_c, x70, x71_c, x72, x74, x76, x77_c, x78_c, x80, x81_c, x82, x83, x84_c, x85_c, x86, x87, x88, x89, x90_c, x92, x94, x95_c, x96_c, x99);
and (w440, x0, x2, x3, x4_c, x5, x6_c, x7, x8, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16_c, x17, x18, x19_c, x20, x21_c, x22_c, x24_c, x25, x26, x27, x28, x30_c, x31, x32_c, x33_c, x34, x36, x37_c, x38, x40_c, x41, x42_c, x43_c, x45, x47_c, x48, x49, x50, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x57_c, x58, x59, x60_c, x61, x62, x63, x64_c, x66, x67, x69, x70_c, x71, x72_c, x74, x75, x76_c, x77_c, x78_c, x79, x80, x81, x82_c, x83_c, x84_c, x86, x87_c, x88_c, x89_c, x90, x91, x92_c, x93_c, x94_c, x95_c, x96, x97, x98, x99);
and (w441, x2_c, x3_c, x4, x5, x7_c, x8, x9_c, x10, x11_c, x12_c, x14, x15, x16, x17, x18, x20_c, x21_c, x23_c, x24_c, x25_c, x26, x27_c, x28, x29_c, x30, x32, x33_c, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x42_c, x43, x44_c, x46, x47_c, x48, x49, x50, x53, x54, x55, x56_c, x57_c, x59_c, x60_c, x63_c, x64_c, x65_c, x66, x67, x68, x69, x70_c, x71_c, x73_c, x75_c, x76, x77_c, x78, x79, x80_c, x81_c, x82_c, x83, x84, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94, x95_c, x96, x97, x98);
and (w442, x0, x1, x2, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x16, x17, x18_c, x20, x21_c, x22, x23_c, x24_c, x25, x27_c, x28, x31_c, x32, x33, x35, x38_c, x39_c, x41_c, x42_c, x43_c, x44, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53, x54, x55, x56, x58, x60, x61_c, x62_c, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x82, x83, x85_c, x87_c, x88_c, x89, x90_c, x91, x92_c, x93_c, x96_c, x97, x98, x99_c);
and (w443, x15, x17_c, x25_c, x27, x32_c, x33_c, x34, x38, x40_c, x42_c, x43_c, x44_c, x66_c, x68, x74_c, x75, x89_c, x97_c);
and (w444, x1_c, x9, x11, x14, x16, x22_c, x25_c, x35_c, x48_c, x55_c, x63_c, x64, x70, x75, x80_c, x85_c, x90_c, x92_c, x96_c, x97);
and (w445, x0_c, x2_c, x3, x5_c, x6, x7, x9, x10_c, x11, x13, x14_c, x15, x16, x17, x18, x19, x21, x22, x25_c, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x35, x37_c, x39_c, x40, x42_c, x43, x44, x45_c, x47, x48_c, x49_c, x50_c, x51, x53, x54_c, x55_c, x56_c, x57, x58, x60, x61, x62_c, x63_c, x64_c, x65_c, x67_c, x68, x69, x70, x71_c, x72, x73_c, x75_c, x76, x77_c, x79_c, x81, x83, x84, x85_c, x87_c, x88, x90, x92_c, x93_c, x94, x95, x96_c, x99_c);
and (w446, x0_c, x1, x2_c, x3, x5_c, x7, x8_c, x9_c, x12, x13_c, x16_c, x17, x18, x19, x20_c, x21_c, x23, x24_c, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x33_c, x34, x35, x36, x37, x38, x40, x41, x44_c, x45_c, x46, x49, x50, x51_c, x52, x53_c, x54_c, x55, x56, x57_c, x58, x60, x63_c, x65_c, x66, x69, x70_c, x71_c, x74_c, x75, x76_c, x77_c, x80, x81, x82_c, x84_c, x85, x86, x87, x90, x93, x94_c, x96, x97);
and (w447, x10_c, x16_c, x19, x29_c, x31, x33_c, x34, x42_c, x48_c, x54_c, x60_c, x64_c, x75_c, x85, x88_c, x89, x98, x99);
and (w448, x1, x2, x3, x4_c, x8_c, x9, x13_c, x14, x17, x18, x19_c, x20_c, x21, x24, x26, x28, x29_c, x30_c, x31_c, x32_c, x33, x34, x37, x38_c, x40, x41, x43_c, x47, x48_c, x49, x51, x52_c, x54_c, x55, x56_c, x59_c, x60, x61_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x70, x72, x73, x75, x77, x78, x79, x80_c, x81, x82_c, x84_c, x87, x89_c, x90_c, x91, x92, x93_c, x94_c, x95, x98, x99);
and (w449, x0_c, x1_c, x2_c, x10_c, x12, x13_c, x20, x21_c, x22_c, x23_c, x26_c, x28_c, x29, x30, x37, x38_c, x39_c, x41, x44_c, x45_c, x50, x51_c, x52_c, x55, x56_c, x59, x61_c, x62, x63_c, x64_c, x65_c, x68_c, x71_c, x72, x74, x78, x80_c, x82, x83_c, x84, x86_c, x87_c, x91, x99);
and (w450, x3_c, x8_c, x12, x14_c, x15_c, x18, x19, x21, x22, x23, x24, x25, x28, x31, x32, x34, x37_c, x41_c, x43_c, x44_c, x46, x50, x51, x52, x53, x54_c, x55_c, x56, x57, x62_c, x63, x64, x68, x71_c, x73_c, x78_c, x79, x80, x81_c, x85_c, x88_c, x90_c, x91, x92, x95, x97_c);
and (w451, x0_c, x1, x2_c, x3_c, x5, x7_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16_c, x17_c, x18, x19, x20, x21, x22_c, x23, x24, x25, x26, x27_c, x28_c, x29, x31_c, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39, x40_c, x41, x42, x43, x44_c, x45, x46, x47_c, x49_c, x50, x51_c, x52_c, x53, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x67, x68_c, x69_c, x70_c, x71_c, x72_c, x73, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83, x84_c, x86, x87, x88, x89_c, x90_c, x91, x92_c, x93, x94, x95, x96_c, x97, x98, x99_c);
and (w452, x0_c, x3, x4_c, x5, x6, x7, x8, x10_c, x11_c, x12_c, x13, x14, x17, x20_c, x22_c, x24_c, x27_c, x28_c, x29, x30_c, x31_c, x32, x38_c, x39, x40, x41, x42, x44, x45_c, x46_c, x50, x51_c, x55_c, x57, x59, x63, x70_c, x71, x72_c, x74_c, x75, x76, x77_c, x80_c, x82, x85, x86_c, x87, x88, x89, x90, x93, x94, x96, x97_c);
and (w453, x0_c, x4, x8_c, x10, x12, x23_c, x27_c, x37_c, x39, x43_c, x46_c, x67_c, x69, x76, x81, x82_c, x84_c, x92, x95);
and (w454, x0, x1_c, x2, x3, x4, x5, x6, x7, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22, x23, x24, x25, x26_c, x27_c, x28, x29, x30_c, x31, x32, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40, x41, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62, x63_c, x64, x65, x66, x67_c, x68_c, x69_c, x70, x71_c, x72_c, x73, x74_c, x75_c, x76_c, x78, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95_c, x96, x97, x98, x99);
and (w455, x1, x2_c, x5, x7_c, x8, x9_c, x10_c, x12_c, x13, x16, x17_c, x18_c, x19, x20_c, x21, x22_c, x23_c, x24_c, x25, x26_c, x27_c, x28_c, x30_c, x31_c, x32_c, x38_c, x40_c, x41, x42_c, x44_c, x45_c, x48, x51_c, x52_c, x53_c, x54, x55, x56, x61, x62_c, x63_c, x64, x65, x66, x68, x69, x72, x73, x74, x75_c, x78, x80_c, x81, x82_c, x84, x85_c, x87, x88, x89, x90_c, x91, x92_c, x93, x97, x99);
and (w456, x26_c, x58_c, x62_c, x70, x94);
and (w457, x1, x2, x5, x6_c, x7_c, x8, x9_c, x10_c, x11, x12, x13_c, x14, x16_c, x18, x20, x21, x22_c, x24_c, x26, x27, x30_c, x31, x32, x33, x35, x37_c, x38_c, x40_c, x42, x43_c, x46_c, x47, x48_c, x49_c, x52_c, x55_c, x57, x59, x60_c, x61_c, x62_c, x63, x64_c, x66, x67, x68_c, x69, x72_c, x73, x75_c, x78, x79, x80, x82_c, x83_c, x84, x86, x87_c, x91, x93, x94, x95, x96_c, x97, x98_c, x99);
and (w458, x1, x4_c, x6, x8, x11_c, x12_c, x15_c, x17, x20_c, x21_c, x24, x27_c, x28, x37, x39_c, x41_c, x43_c, x47, x49, x50, x52_c, x53_c, x57_c, x62_c, x69_c, x73, x76_c, x81, x82_c, x86, x88_c, x89_c, x90, x91_c, x93, x94, x95);
and (w459, x1_c, x2, x4, x5_c, x6_c, x8_c, x11, x12_c, x16_c, x17_c, x18, x19, x21, x22_c, x23_c, x24_c, x27_c, x29, x31, x32_c, x33_c, x34, x35, x36_c, x37_c, x40_c, x42_c, x44_c, x45, x47, x49, x50, x53, x54, x55_c, x56, x57_c, x59, x61, x62, x64_c, x65, x69, x70_c, x71_c, x72, x73_c, x74, x75_c, x79_c, x80, x81_c, x82_c, x85_c, x86_c, x89_c, x91, x92_c, x94_c, x96_c, x97_c, x98_c, x99_c);
and (w460, x6_c, x8, x12_c, x17_c, x24_c, x26_c, x36, x37_c, x42_c, x43, x48, x49_c, x51, x71, x73_c, x75_c, x76, x80, x95_c, x99);
and (w461, x0_c, x1, x2, x3_c, x4_c, x5, x6, x7, x8, x9, x10, x11_c, x12, x13, x15, x16, x17_c, x18_c, x19, x20_c, x22, x24, x25_c, x26_c, x27_c, x28, x29_c, x30, x31, x32_c, x33, x34, x35, x36_c, x37, x38_c, x40_c, x41, x42, x43, x44_c, x45_c, x46, x47_c, x48, x49, x50_c, x51, x52_c, x53_c, x54_c, x55_c, x57, x59_c, x60, x61_c, x62, x63, x64, x65_c, x66, x67_c, x68_c, x69, x70_c, x71_c, x72, x73_c, x74_c, x75_c, x77, x78, x79_c, x81, x82, x83_c, x84_c, x85_c, x86, x88, x89_c, x90, x91_c, x92_c, x93, x94_c, x96, x97_c, x98, x99);
and (w462, x0_c, x3_c, x4_c, x6, x7_c, x10, x11, x13, x16, x17_c, x18, x20_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31_c, x33_c, x35, x36, x40, x41_c, x42, x43_c, x44_c, x45, x47, x48, x50, x52_c, x53_c, x54, x55_c, x56_c, x60, x63_c, x64, x65_c, x67_c, x70, x73_c, x74_c, x77_c, x81_c, x82, x83_c, x85_c, x86_c, x87_c, x88, x91_c, x92, x93, x94_c, x96, x98);
and (w463, x0, x2_c, x5_c, x9, x10, x13, x15, x18, x22, x26_c, x29, x30, x31, x33, x35_c, x39, x40_c, x41, x42, x45, x46, x48_c, x49_c, x52_c, x57_c, x59, x60, x62_c, x63_c, x66, x69, x70_c, x72, x73, x74_c, x75, x79, x81, x87, x90, x91, x92, x93, x94_c, x96_c);
and (w464, x0_c, x1_c, x3_c, x5_c, x7_c, x10, x11_c, x14, x19_c, x21, x23, x24_c, x29, x30, x31, x34, x36, x39_c, x40, x41, x44_c, x46_c, x47, x49_c, x50_c, x59, x63_c, x66, x68_c, x70_c, x73_c, x75_c, x77_c, x78, x79, x80_c, x81, x83_c, x84, x86_c, x88, x90_c, x93_c, x94_c, x96, x97, x98);
and (w465, x2_c, x6, x8_c, x12_c, x13_c, x15_c, x16_c, x18_c, x24, x26_c, x31_c, x34, x35_c, x52_c, x56_c, x62, x64, x69, x75, x77, x88_c, x89_c, x95);
and (w466, x0, x1_c, x2_c, x3, x4, x5, x6, x7_c, x8_c, x9_c, x10, x12_c, x13_c, x15_c, x16, x18_c, x19, x21, x23_c, x24, x25, x26, x27, x28_c, x30_c, x31_c, x32, x33, x34_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x45_c, x47_c, x48, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x57_c, x58_c, x60_c, x61, x62, x63_c, x65_c, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75, x76, x77_c, x78_c, x80, x82, x83_c, x84, x85, x86_c, x87, x88_c, x90_c, x91_c, x92_c, x93_c, x94_c, x97, x98, x99_c);
and (w467, x7, x9_c, x11, x12_c, x13_c, x17, x26, x27, x29_c, x30, x32, x36_c, x40_c, x41_c, x42, x43, x46, x47, x48_c, x49_c, x52_c, x53, x57, x58_c, x60, x61, x62, x63_c, x64_c, x65, x67, x68_c, x70, x71, x72_c, x73, x74, x77_c, x82_c, x83_c, x86_c, x87, x88, x89, x90_c, x92, x93_c, x94_c, x96, x97_c, x99);
and (w468, x31_c, x36, x38_c, x47, x63, x67_c, x69_c, x75_c, x89);
and (w469, x3_c, x18, x27_c, x34_c, x73_c, x98);
and (w470, x2_c, x3_c, x6, x10, x11, x19, x20_c, x22, x24, x25, x26, x28, x31_c, x33, x34_c, x37, x38_c, x39, x43_c, x45, x46, x50_c, x61, x67, x70_c, x73, x74_c, x76, x81_c, x85, x89, x92_c, x95, x97, x98_c);
and (w471, x6_c, x8, x17_c, x26_c, x37, x44, x47_c, x62, x69);
and (w472, x1, x7, x20_c, x24, x25, x29_c, x44, x56, x71, x91_c, x94, x96_c, x98_c);
and (w473, x8, x17, x18_c, x27_c, x34, x39_c, x55, x56_c, x61_c, x62_c, x70_c, x88_c);
and (w474, x0_c, x1, x2, x3_c, x4_c, x5_c, x6, x7, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15, x16_c, x17, x18, x19_c, x20, x21_c, x22_c, x23, x24, x25, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x42_c, x43, x45_c, x46_c, x47, x48_c, x50_c, x51, x52_c, x53_c, x54, x55, x56_c, x57_c, x58_c, x59_c, x60, x61, x62_c, x63_c, x64, x66, x67_c, x68_c, x69_c, x70_c, x71_c, x72, x73, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81_c, x82, x83, x84, x85, x86, x87_c, x88, x90_c, x91, x92_c, x93_c, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w475, x2_c, x3_c, x4, x5, x6_c, x8, x9_c, x11_c, x12_c, x13, x14_c, x19_c, x21_c, x24_c, x28, x30, x31, x32, x35_c, x36, x39_c, x40_c, x41_c, x42, x43, x44_c, x45_c, x46, x48, x51_c, x52_c, x53, x54, x55, x57, x60_c, x61_c, x62, x63, x65_c, x68, x69, x72_c, x73, x76, x78, x79_c, x81, x82, x84_c, x86_c, x87, x90, x94, x95, x96, x97, x98);
and (w476, x2, x3_c, x9, x13, x14, x15, x20, x35, x37, x38_c, x39_c, x40_c, x41_c, x43_c, x44_c, x45_c, x46_c, x47_c, x51, x53, x55, x57_c, x59, x61, x64_c, x65, x66_c, x72_c, x76_c, x82_c, x84_c, x85, x86, x88_c, x92_c, x93);
and (w477, x0, x1, x2, x3_c, x4, x5, x6_c, x7, x8_c, x9, x12, x13, x15, x16, x18_c, x19_c, x20, x22, x23_c, x24, x26_c, x27_c, x28_c, x29_c, x30, x32, x34, x35_c, x36_c, x37, x38_c, x40, x42, x43, x44, x45_c, x46_c, x47_c, x48, x50_c, x51_c, x56, x57_c, x59_c, x60_c, x61, x62, x63_c, x64, x66_c, x67, x70_c, x72, x74_c, x75, x77, x78, x80_c, x81, x82, x83, x86, x88, x89_c, x91, x92, x93, x94_c, x95, x96_c, x97_c, x99_c);
and (w478, x0_c, x1_c, x2_c, x4_c, x5, x6, x7_c, x9, x13, x14_c, x16_c, x17, x18, x20_c, x22_c, x23, x24_c, x25, x26_c, x28, x29_c, x31_c, x32_c, x35_c, x37, x38, x40_c, x41_c, x43_c, x47, x49, x50_c, x52_c, x53_c, x54, x55_c, x56, x58, x59_c, x60, x62, x63, x64, x66, x68, x69_c, x70, x71, x72, x74_c, x75_c, x76_c, x77_c, x78, x82, x85, x88, x89, x90_c, x91, x92_c, x93_c, x94_c, x95, x98_c, x99_c);
and (w479, x6, x17_c, x20_c, x24_c, x25_c, x27_c, x28_c, x32, x41_c, x44, x50, x52_c, x57_c, x61_c, x62, x64, x65, x69, x77, x81, x88, x89, x90_c, x92_c, x94, x95_c);
and (w480, x8, x30_c, x38, x41_c, x49, x56_c, x87, x92_c);
and (w481, x60_c, x69_c);
and (w482, x3, x4_c, x6_c, x12_c, x16_c, x23_c, x24_c, x29_c, x31_c, x36_c, x39_c, x45_c, x46, x50_c, x53, x54, x55_c, x56, x62, x68, x70_c, x72_c, x81_c, x83, x89_c, x91, x92_c, x93_c, x96, x97_c);
and (w483, x3_c, x7_c, x9_c, x12_c, x15, x17, x18_c, x22, x24_c, x27_c, x30, x32, x33_c, x34_c, x35_c, x37_c, x39_c, x40_c, x41_c, x45_c, x46_c, x47, x49, x52_c, x54_c, x55, x56_c, x58, x59_c, x60_c, x61, x62, x64_c, x66, x68, x72_c, x73, x74_c, x76, x77, x80, x81, x86_c, x88, x90, x92, x95_c, x96);
and (w484, x0_c, x1_c, x2, x3, x8, x9_c, x12_c, x13_c, x14_c, x15_c, x18_c, x19, x20_c, x24_c, x26_c, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x35, x37_c, x38_c, x39, x41, x44, x45_c, x46_c, x48, x49_c, x52, x53, x60_c, x62_c, x63, x67_c, x70, x71, x74_c, x75, x76, x78_c, x80_c, x83_c, x84, x86, x88_c, x93_c, x95);
and (w485, x2_c, x3, x4, x6_c, x11, x12, x13, x15, x16_c, x20_c, x22, x23, x24_c, x25, x32_c, x33_c, x34_c, x38, x39_c, x43_c, x45, x46_c, x49_c, x50, x56, x57_c, x58, x59, x62_c, x64_c, x66, x67_c, x70_c, x73, x74_c, x79, x80, x83_c, x84, x85_c, x86, x90_c, x91, x93_c, x94);
and (w486, x3_c, x4, x5, x8, x10, x13, x15_c, x17_c, x18, x19_c, x20_c, x21, x23, x24, x25, x27, x30_c, x31, x37_c, x42_c, x44_c, x45_c, x47_c, x49_c, x50_c, x54_c, x55, x58_c, x60, x61_c, x64, x66, x69, x70, x73, x75, x76, x77, x80_c, x81, x83, x86_c, x91, x92, x96, x98, x99);
and (w487, x2_c, x8_c, x15_c, x26, x35, x36, x51, x54_c, x69_c, x70, x71, x77, x79, x82_c, x84_c, x93_c, x94, x95, x96_c, x98);
and (w488, x0, x1_c, x2_c, x3_c, x4, x5, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x14, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23_c, x25, x26, x27, x28_c, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39, x40, x42, x43, x44_c, x45_c, x46_c, x47, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62_c, x65_c, x66_c, x67, x68_c, x70, x71, x72_c, x73, x74, x75, x76_c, x77_c, x79_c, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88, x89_c, x90, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w489, x20_c, x25_c, x32, x53, x55_c, x57_c, x77_c, x79_c);
and (w490, x9_c, x17_c, x26, x27, x28_c, x33_c, x34, x39, x47_c, x49_c, x51, x56_c, x59, x62_c, x68, x99_c);
and (w491, x2, x6_c, x7_c, x8, x10, x12_c, x13, x14_c, x15, x17, x19_c, x20_c, x22, x23_c, x24, x25, x29, x30, x34, x36, x40_c, x42_c, x50_c, x51, x52, x55_c, x56_c, x57, x58, x59_c, x60_c, x61, x62_c, x65, x66, x67, x69, x75, x79, x80_c, x81_c, x82_c, x89, x91, x92, x95_c, x96, x97);
and (w492, x0, x5, x6_c, x7, x9_c, x10_c, x12_c, x14, x15_c, x16_c, x17_c, x18, x20, x21, x22, x25, x26_c, x27_c, x29, x30_c, x32_c, x33, x34_c, x36, x37_c, x38, x39, x40, x42_c, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50, x52_c, x53, x54, x55_c, x56_c, x57, x59, x60_c, x61_c, x63_c, x64_c, x65_c, x66, x67, x68, x69_c, x70, x71_c, x74_c, x75_c, x76, x77, x78, x79, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86, x87_c, x88, x89, x91, x92, x95_c, x96_c, x98_c, x99);
and (w493, x0, x2_c, x3, x4_c, x5_c, x8_c, x10, x11, x15_c, x18, x29, x33, x40, x41_c, x47_c, x51, x52_c, x53_c, x56_c, x57, x61, x63_c, x64, x67, x69, x70_c, x73_c, x83, x84, x86_c, x87_c, x88_c, x90, x93_c, x94, x95, x97_c, x98, x99);
and (w494, x3, x4_c, x9, x15_c, x16_c, x19_c, x20_c, x21_c, x22_c, x24, x27_c, x33, x37_c, x43_c, x44, x58_c, x63_c, x67, x72_c, x77_c, x80_c, x84, x90_c, x93, x99);
and (w495, x1_c, x2, x7, x13, x19_c, x20_c, x23_c, x24_c, x29_c, x35, x39_c, x45_c, x54, x61_c, x69, x70_c, x71_c, x73_c, x79, x81, x85_c, x90, x92, x97, x99_c);
and (w496, x1, x2_c, x3_c, x6_c, x7, x8, x9_c, x10, x11_c, x12, x15_c, x16, x17, x18_c, x22, x25_c, x26, x34, x35_c, x36_c, x37, x39, x40, x41_c, x42, x47, x48, x49, x51_c, x61_c, x68_c, x69, x71, x72, x74_c, x75, x78_c, x79_c, x88_c, x91_c, x92_c, x93, x94, x95, x96, x97, x98_c, x99);
and (w497, x5, x9_c, x11_c, x12_c, x14, x18, x20, x26, x30, x32, x33, x35, x42, x44, x45, x47, x48_c, x51_c, x53_c, x55_c, x58, x59, x66_c, x70, x71_c, x73_c, x74_c, x75_c, x80_c, x82, x83_c, x86_c, x94, x98_c);
and (w498, x0, x3_c, x4, x5_c, x6_c, x8_c, x13, x20_c, x28_c, x37_c, x38, x41, x43_c, x44, x45_c, x47_c, x50, x56_c, x58_c, x60, x61, x62, x63, x66_c, x67_c, x72_c, x73, x75, x78_c, x81_c, x85, x87, x88, x97_c);
and (w499, x10, x13_c, x14, x30, x33_c, x34_c, x42_c, x45, x51, x56_c, x64, x68, x71_c, x72_c, x73_c, x75_c, x77, x79, x80_c, x94);
and (w500, x3_c, x4, x7, x9_c, x23, x25, x26_c, x28_c, x30, x44_c, x49, x50_c, x52, x53, x54, x57_c, x61_c, x65_c, x68, x70, x73, x78, x80_c, x81, x82_c, x83, x89, x90_c, x92, x93_c, x95, x96_c);
and (w501, x0_c, x2, x4_c, x7, x10, x15, x16_c, x20_c, x22_c, x23_c, x29, x30, x31_c, x37_c, x41, x44_c, x48_c, x51_c, x52, x54_c, x55, x56, x57, x61_c, x62, x65, x70, x73, x74, x75_c, x78, x79_c, x81, x85, x88, x91_c, x93, x99_c);
and (w502, x0_c, x1_c, x2, x3_c, x4, x6, x7_c, x8, x9, x10_c, x12_c, x13_c, x14, x15, x16, x17_c, x18, x19, x20, x21, x23, x24_c, x25_c, x26_c, x28_c, x29_c, x30, x32, x33, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42, x43_c, x44_c, x45_c, x47_c, x48_c, x50, x51, x52, x53, x54, x55, x56_c, x57_c, x58, x59_c, x60, x61_c, x62_c, x63, x64_c, x65, x66, x68, x69, x70, x71, x72_c, x73, x74_c, x75_c, x76_c, x77, x78_c, x79, x80, x81, x82, x83, x84_c, x86, x87_c, x88_c, x89, x90_c, x91, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w503, x1_c, x2, x3, x5_c, x6, x8_c, x9, x11_c, x12_c, x13_c, x17, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35_c, x36, x37, x38, x40_c, x42_c, x47_c, x48, x49, x54_c, x56_c, x59, x63, x64_c, x67, x68, x69_c, x70_c, x73_c, x74_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84, x86_c, x87_c, x90, x92, x94, x95, x96_c, x97, x98);
and (w504, x0, x1_c, x2, x3_c, x4, x5_c, x6, x7_c, x9_c, x10_c, x14, x15, x16, x17, x18_c, x19, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27_c, x28, x29, x31_c, x32_c, x34_c, x35_c, x36, x38, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x47_c, x48, x49_c, x51, x52_c, x54_c, x55, x57, x58_c, x59_c, x60, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69, x70, x71_c, x73, x74, x75, x76, x77_c, x78, x79_c, x80, x81_c, x82_c, x83, x84_c, x85_c, x87_c, x88_c, x90_c, x91, x93, x95, x96, x97, x98_c, x99);
and (w505, x0_c, x1, x2_c, x4, x7, x9_c, x12_c, x13, x15_c, x16, x17, x18, x19_c, x20_c, x21_c, x22_c, x23, x26_c, x28, x31, x32, x34, x36, x39_c, x40, x41, x42_c, x44_c, x45_c, x46_c, x49_c, x50_c, x51_c, x52, x53, x54, x55, x57_c, x58_c, x61_c, x62, x63, x64, x65_c, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x73, x76_c, x77_c, x81_c, x82, x83, x86, x88, x89, x90, x91_c, x93, x94, x95_c, x96_c, x97, x98, x99);
and (w506, x4, x38_c, x41, x78_c, x85);
and (w507, x0_c, x1_c, x2, x3_c, x6, x8, x9, x10, x11, x12, x13, x15, x16, x18_c, x20_c, x21, x22_c, x23, x26, x28, x31_c, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x40, x43_c, x44, x45_c, x49_c, x52, x53_c, x55, x57, x58, x60, x61, x63_c, x66, x68_c, x70, x71, x74, x75, x76_c, x77, x79_c, x81, x82, x84, x85, x86_c, x88, x89_c, x91_c, x92, x93_c, x94, x95_c, x96, x98);
and (w508, x2, x3_c, x4_c, x6_c, x7_c, x8_c, x10, x14, x15, x16, x18, x20, x21, x22_c, x25_c, x29, x31_c, x32_c, x33, x34_c, x35_c, x39_c, x41_c, x42_c, x44, x45_c, x46, x47, x48, x49, x50_c, x51_c, x52_c, x54, x55_c, x56_c, x58, x59, x60, x61_c, x62_c, x64_c, x67_c, x69_c, x73_c, x76_c, x78_c, x84, x86, x90_c, x91_c, x95, x96, x98_c);
and (w509, x1, x3_c, x4_c, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12, x13_c, x16, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x28_c, x29_c, x30, x31, x32, x33, x39, x40, x42_c, x44, x45_c, x46_c, x47, x48, x49, x50, x51, x52_c, x54_c, x55, x56_c, x57_c, x58_c, x60_c, x61_c, x62, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x69, x70, x71, x73_c, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83, x84_c, x85, x86_c, x87, x88, x89, x90_c, x91, x92_c, x93, x94, x95_c, x96_c, x97_c, x98, x99_c);
and (w510, x51_c, x58_c, x65);
and (w511, x1, x7, x9, x10_c, x11, x13_c, x14, x15, x17_c, x19, x20_c, x22, x25, x27_c, x29_c, x31_c, x32, x33, x34_c, x39, x40, x43_c, x45, x48, x52_c, x60_c, x61, x67_c, x68_c, x69_c, x70_c, x71_c, x72_c, x76_c, x78, x79, x82, x83, x84_c, x85, x89_c, x97, x98);
and (w512, x0_c, x2, x3, x4, x5_c, x9_c, x12_c, x13, x15_c, x16_c, x17_c, x18_c, x21, x22, x23, x25_c, x27, x28, x29, x30_c, x33_c, x34_c, x35, x39_c, x41, x43, x45_c, x46_c, x47, x50_c, x52, x53, x54_c, x55, x61_c, x63, x64_c, x65_c, x67, x68, x69, x71_c, x72, x76_c, x77_c, x79, x81, x82, x83, x84_c, x88, x89, x91, x92_c, x95_c, x96, x97, x98, x99);
and (w513, x0, x3_c, x13_c, x15, x16_c, x17, x19_c, x23_c, x25, x46_c, x50_c, x54_c, x58_c, x59, x67_c, x72_c, x76_c, x85, x86, x94, x99_c);
and (w514, x0, x1, x2_c, x3, x8_c, x9, x13, x14, x15_c, x16, x17_c, x18_c, x20, x22, x23, x25_c, x28_c, x29_c, x30_c, x31, x34, x35_c, x37_c, x38, x40_c, x42, x44, x45_c, x47, x49_c, x50_c, x53, x56, x58, x59, x60_c, x61_c, x62, x66_c, x67, x68_c, x71_c, x73_c, x74, x75_c, x76_c, x77, x79, x81_c, x82_c, x83_c, x84_c, x85_c, x87, x91_c, x92, x94, x95, x96_c, x98_c, x99);
and (w515, x0, x1_c, x3, x4_c, x6, x7_c, x8_c, x9_c, x10, x11_c, x12, x13, x14, x15_c, x16, x17_c, x18, x20_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x30, x33, x34_c, x35_c, x38, x43_c, x44, x45, x47, x48, x49, x50_c, x51, x52_c, x53, x54, x55, x58_c, x59, x61, x62_c, x64, x65_c, x67, x69_c, x70_c, x71_c, x73, x74_c, x75_c, x76, x79, x80, x81, x82, x85_c, x86_c, x87_c, x88, x90, x91_c, x92_c, x93_c, x94_c, x95, x97, x98, x99);
and (w516, x0, x1_c, x2_c, x3, x4_c, x5, x7, x8_c, x10, x12, x13_c, x14, x16_c, x17, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x33, x34_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x43, x44, x45_c, x46_c, x47, x48, x49_c, x50, x51_c, x52_c, x53, x54_c, x55, x56_c, x57, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x67, x68_c, x70_c, x71, x72, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79, x80_c, x81_c, x82, x83, x84, x85, x86_c, x88, x89, x90_c, x91, x92_c, x93, x94_c, x95, x96_c, x97, x98, x99);
and (w517, x0_c, x1_c, x5_c, x6, x7, x8, x10_c, x11_c, x12, x13_c, x17, x18, x19, x20, x21_c, x26, x27, x30, x31, x32, x33, x35_c, x36, x37, x38_c, x39_c, x40_c, x41, x43_c, x44, x46, x48, x49, x50, x51, x52, x55, x56_c, x57, x58_c, x60, x62, x63, x64_c, x65, x66, x67, x69, x70_c, x71, x72_c, x73, x76, x78_c, x81, x82, x83_c, x84_c, x85, x86, x87_c, x88_c, x90_c, x91, x92_c, x94_c, x95, x96, x97);
and (w518, x0, x1_c, x4_c, x7, x17_c, x18_c, x52_c, x66_c, x67_c, x70_c, x74_c, x99_c);
and (w519, x0, x1, x2_c, x3, x5, x6, x7, x8, x9, x10_c, x11, x13, x14_c, x15_c, x16, x17, x18, x20_c, x23, x24_c, x26_c, x28_c, x29_c, x30_c, x31, x32, x33, x35, x36, x37_c, x38_c, x39_c, x40_c, x41, x42_c, x44, x47_c, x48_c, x50, x51, x52, x53_c, x54_c, x55_c, x56, x57_c, x59_c, x61, x62, x64, x65, x66, x68_c, x69, x70_c, x73, x74, x76, x77, x78, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85, x86, x89, x91_c, x92_c, x93_c, x95, x96_c, x97_c, x99_c);
and (w520, x3, x11, x27, x34_c, x40_c);
and (w521, x8, x14_c, x16_c, x18, x22, x23_c, x27_c, x37, x38_c, x40, x51_c, x57, x62, x65_c, x70, x71_c, x72_c, x73_c, x76, x79_c, x83, x90);
and (w522, x7_c, x9_c, x12_c, x14_c, x15_c, x16, x18, x19_c, x20_c, x22, x23_c, x24_c, x25, x30, x31_c, x32_c, x35_c, x36_c, x38_c, x39, x40, x41_c, x44_c, x46_c, x47_c, x48, x49_c, x51_c, x61, x62_c, x63_c, x65_c, x66_c, x68, x69_c, x71, x73, x74, x75_c, x77, x78, x79, x82_c, x84_c, x85, x88, x89, x90, x91, x92_c, x94, x96, x99_c);
and (w523, x0, x6, x7_c, x9, x10, x15_c, x32_c, x36, x51_c, x63, x69_c, x70, x72, x78_c, x89_c, x92_c, x97);
and (w524, x4_c, x33, x44);
and (w525, x0_c, x1, x2_c, x3, x4, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25, x26, x27_c, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36_c, x37_c, x38, x39_c, x40_c, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48, x49, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56_c, x57_c, x58, x59, x60, x61, x62, x63_c, x64_c, x65_c, x66, x67, x68_c, x69, x70_c, x71, x72, x73, x74, x75_c, x76, x77, x78, x79_c, x80_c, x81, x82_c, x83, x84, x85, x86, x87_c, x88_c, x89, x90_c, x92_c, x93_c, x94, x95, x96, x97, x98, x99);
and (w526, x1, x3_c, x4, x5_c, x6_c, x7_c, x9_c, x12_c, x15_c, x16, x17, x18, x19_c, x20_c, x21_c, x27, x29_c, x30_c, x32, x35_c, x39, x40, x42, x44_c, x46, x50, x51_c, x53_c, x55, x56_c, x60, x70_c, x72_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x92_c, x97_c, x99_c);
and (w527, x0_c, x3_c, x5_c, x6, x10, x13_c, x14, x16_c, x17_c, x23_c, x25, x27, x28_c, x29, x31_c, x36, x38_c, x40, x44, x50_c, x51, x55_c, x56_c, x58, x59_c, x61, x62, x63_c, x64_c, x73, x74_c, x75_c, x76_c, x77_c, x79, x81_c, x82, x89, x90_c, x91_c, x93, x94_c, x96, x97_c, x98);
and (w528, x15, x24, x33, x37_c, x56_c, x65_c, x82, x94, x98);
and (w529, x0_c, x2_c, x3_c, x6_c, x7, x8, x9_c, x10, x11_c, x12_c, x13_c, x14, x16_c, x17, x18, x19_c, x22_c, x23_c, x24_c, x27, x28_c, x29, x31, x32_c, x33, x34, x35, x36, x38, x39, x40_c, x41_c, x42, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51_c, x54, x55, x58, x59, x60, x61_c, x63, x64, x65_c, x66_c, x67_c, x69_c, x70, x71, x72, x73_c, x74, x75_c, x77_c, x78, x79, x81_c, x82, x83_c, x84, x85_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99);
and (w530, x0, x1, x2, x3_c, x4, x6, x9, x10_c, x11_c, x12_c, x13_c, x14_c, x17, x19, x20_c, x21_c, x22, x23, x24_c, x25_c, x26_c, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34_c, x35, x36, x37_c, x38, x39, x40_c, x41_c, x43, x44_c, x45_c, x46_c, x47, x48_c, x49, x51_c, x52, x53, x54_c, x55_c, x58, x60_c, x61, x62, x64, x65_c, x67, x68_c, x69_c, x70_c, x71, x72, x74_c, x76_c, x77_c, x78_c, x79, x80_c, x81_c, x82, x83, x84, x85, x86_c, x87, x88_c, x89_c, x91, x92, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w531, x6, x15, x17, x19_c, x40_c, x43, x45_c, x48, x55_c, x58_c, x62_c, x67_c, x78_c, x94);
and (w532, x0_c, x2, x4_c, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x18_c, x19, x21, x22, x25, x26_c, x27, x28, x29, x31, x33_c, x34_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51, x53_c, x54_c, x56_c, x58, x59, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80, x81, x83_c, x85_c, x86_c, x87_c, x90, x91, x92, x93, x94_c, x95, x96_c, x97, x98, x99_c);
and (w533, x0, x1_c, x7, x9, x10_c, x12, x13_c, x14, x16, x19, x20, x21, x22_c, x24, x25_c, x26, x29, x30, x34_c, x35_c, x36_c, x37, x38_c, x41, x43, x48, x50_c, x52, x53_c, x54_c, x55, x56_c, x57_c, x58_c, x61_c, x65_c, x66, x67, x68_c, x69, x70, x72, x73_c, x75_c, x77_c, x78, x79, x83_c, x84, x86_c, x87_c, x89_c, x90_c, x92_c, x93, x94, x95, x98_c);
and (w534, x0_c, x1_c, x2, x3, x4_c, x5, x6_c, x7_c, x8, x9, x10_c, x11_c, x12, x13, x14_c, x15_c, x16, x17_c, x19_c, x20, x21_c, x22, x23_c, x24, x25, x26, x27_c, x29_c, x31_c, x32, x33_c, x35_c, x36, x37, x38, x40, x41_c, x42_c, x43_c, x44, x46_c, x47_c, x48, x50_c, x51, x52, x53, x54, x55, x56, x57, x58_c, x59, x61_c, x62, x63_c, x64, x65, x66_c, x67_c, x68_c, x69_c, x71, x72, x77, x78, x79_c, x80, x81, x82, x83, x84, x87_c, x88, x89_c, x91, x92, x95, x96, x97, x98, x99_c);
and (w535, x0, x1_c, x2, x7_c, x8_c, x10_c, x13_c, x14, x15_c, x16_c, x17_c, x20_c, x21_c, x24, x25_c, x26_c, x28, x30_c, x32, x34, x38_c, x42_c, x43, x50, x53_c, x55, x57_c, x58_c, x59, x61_c, x62_c, x63_c, x64_c, x65, x67, x69_c, x70_c, x72_c, x73_c, x74_c, x77_c, x79_c, x87_c, x92, x94_c, x95_c, x96_c, x97);
and (w536, x1, x5_c, x10, x12_c, x17, x18_c, x19, x26_c, x31, x37, x44, x53, x54_c, x58_c, x62, x63, x65, x68, x72_c, x73, x74, x75, x84_c, x85, x87, x88, x91_c, x94, x95, x96_c);
and (w537, x0, x1_c, x2, x9, x11, x12, x20, x23_c, x27_c, x29, x32, x33, x41, x47, x48_c, x49, x50_c, x51_c, x52, x55, x56, x59_c, x60_c, x61_c, x62, x64_c, x69, x71_c, x73, x74, x77_c, x86_c, x89, x91, x99);
and (w538, x1_c, x2_c, x7, x13_c, x18_c, x26, x27_c, x38, x40_c, x51_c, x54_c, x55_c, x61, x63_c, x64, x70_c, x71, x74_c, x82_c, x89_c, x91, x93, x94, x97);
and (w539, x0_c, x1_c, x2_c, x4, x5_c, x6_c, x7, x8, x9, x10_c, x11, x12, x13_c, x15_c, x16_c, x19_c, x21_c, x23, x24, x27, x28_c, x30_c, x32, x33_c, x34, x36_c, x37, x38, x39, x41, x42, x45_c, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x54, x55, x57, x58_c, x59_c, x60, x61_c, x62, x63_c, x64_c, x65, x66, x67, x68, x69_c, x70, x73, x75_c, x76_c, x77_c, x78, x79_c, x80, x81_c, x82, x84_c, x85, x86, x87, x89_c, x90, x91_c, x93_c, x94, x95_c, x97, x98, x99_c);
and (w540, x3_c, x5, x7, x8_c, x14, x15_c, x17_c, x21_c, x27_c, x31, x35, x38_c, x39_c, x41, x44_c, x45_c, x47_c, x51_c, x55_c, x58_c, x59_c, x64_c, x66_c, x67_c, x69_c, x76_c, x81_c, x82_c, x85, x99);
and (w541, x1, x8_c, x13_c, x14, x15_c, x16_c, x17, x18_c, x20, x22, x23_c, x24_c, x25_c, x26_c, x27, x29, x30, x32_c, x33, x34, x36, x37_c, x38, x40_c, x54, x58_c, x59_c, x60, x61, x62_c, x63, x64_c, x65_c, x66, x68_c, x69, x70, x71, x73, x76_c, x77, x79, x81_c, x82, x83_c, x84, x85, x90, x92, x93_c, x96, x99_c);
assign w542 = x20_c;
and (w543, x2_c, x5_c, x6_c, x7, x8, x9_c, x10, x11, x12, x13_c, x16, x17, x18, x19_c, x24, x26_c, x27, x29, x31, x33_c, x36, x39_c, x40, x41_c, x42, x43, x44, x45_c, x46, x48_c, x49, x52_c, x53_c, x54_c, x56_c, x57_c, x59_c, x62_c, x64_c, x66_c, x67_c, x68, x72, x75_c, x78, x79, x82, x84, x85_c, x87_c, x88, x89_c, x90_c, x91_c, x92, x93, x95, x96, x97_c, x98_c);
and (w544, x0_c, x1, x2, x3, x4, x5_c, x6, x7_c, x8, x9, x10, x11_c, x12, x14, x16_c, x17, x18, x19, x20, x21, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29_c, x30, x31, x32, x33, x34_c, x36_c, x37, x38_c, x39, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48_c, x49, x50_c, x51_c, x52_c, x53, x54, x55, x56, x57_c, x59, x60, x62_c, x63, x64_c, x65, x66, x67_c, x68, x69, x70_c, x71, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x79_c, x80_c, x81, x82, x83, x84, x85, x86_c, x87, x88, x89_c, x90, x91, x92, x93, x94, x95, x96_c, x97, x98_c, x99_c);
and (w545, x0, x1_c, x3, x4_c, x5, x9_c, x12, x16_c, x18, x20_c, x21, x22, x23, x25, x26_c, x27, x28, x32, x36, x37_c, x38, x40, x45, x48_c, x49, x50_c, x51_c, x55, x56, x57_c, x59, x60, x67, x68_c, x69_c, x71, x72_c, x77_c, x78, x80, x81_c, x82_c, x83, x85_c, x87_c, x88, x90, x91_c, x93, x94_c, x98, x99);
and (w546, x3_c, x11, x15_c, x19_c, x20_c, x21, x24_c, x25, x26_c, x31, x33_c, x34, x36, x44, x49, x57, x62, x64_c, x65, x72, x73, x76_c, x78_c, x85, x88, x89_c, x91_c, x93);
and (w547, x11_c, x15_c, x16, x18, x21, x28_c, x35_c, x36, x37_c, x39, x40_c, x41, x42_c, x44_c, x47_c, x52, x61, x64_c, x65_c, x67_c, x69_c, x70_c, x73_c, x75_c, x79, x80_c, x82, x83_c, x84_c, x91_c, x92);
and (w548, x0_c, x1_c, x2, x3_c, x4, x5, x7, x8_c, x10, x11, x12_c, x13_c, x16_c, x17_c, x19_c, x20_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x28_c, x29, x30, x31, x32, x33_c, x34_c, x35, x36_c, x37_c, x38, x40, x41_c, x43, x44_c, x45_c, x47_c, x48_c, x50_c, x51_c, x53, x54_c, x55_c, x57_c, x58, x59, x61_c, x62_c, x63, x64, x65, x66, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75, x76_c, x77, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84, x85, x86_c, x87, x89, x90, x92, x93, x94, x95, x96_c, x97, x98, x99);
and (w549, x8, x21_c, x25_c, x27_c, x34, x39_c, x44_c, x57, x72, x76_c, x86_c, x88_c, x91, x99);
and (w550, x8_c, x21_c, x44_c);
and (w551, x6_c, x7_c, x8_c, x9, x10, x14_c, x15_c, x20, x21, x22, x26_c, x27, x28, x29_c, x30, x31_c, x32_c, x35_c, x37_c, x38_c, x40_c, x41_c, x42_c, x43_c, x47_c, x48, x51, x53_c, x54, x56, x57_c, x60, x64_c, x65_c, x66, x71_c, x73, x74_c, x75, x77_c, x79_c, x80, x81, x82, x84_c, x86_c, x87_c, x88, x89_c, x92_c, x93_c, x94_c, x95_c, x96_c, x99);
and (w552, x8, x9_c, x16, x24, x25, x26, x32_c, x40, x42_c, x45, x48, x60_c, x63, x69_c, x87, x91, x94, x98_c, x99_c);
and (w553, x0, x1_c, x2_c, x3, x4_c, x5_c, x6, x8_c, x9_c, x10_c, x11, x12, x14, x15, x16, x17_c, x18_c, x19, x20_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x30, x31_c, x32_c, x33_c, x34, x36_c, x37_c, x38_c, x40_c, x41, x42_c, x43, x44_c, x45, x46, x47_c, x48, x49, x50_c, x51_c, x52_c, x53_c, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62, x64, x65_c, x66_c, x67, x68_c, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x75, x77, x78, x79, x80, x81_c, x82_c, x83, x84, x85_c, x86_c, x87, x88, x89, x90_c, x91, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w554, x0_c, x5_c, x6, x12_c, x16, x17_c, x20_c, x21_c, x25_c, x28, x30, x31, x33, x34_c, x38_c, x40, x43, x49, x50, x51_c, x53, x58_c, x61_c, x70_c, x73_c, x85_c, x90_c, x91, x96, x97, x98_c);
and (w555, x1, x3_c, x9, x11_c, x12, x16, x17, x20_c, x21_c, x22_c, x30, x31_c, x32, x33, x44, x47_c, x49_c, x56, x60, x61_c, x65, x66_c, x75_c, x77, x82, x83, x93_c, x97_c);
and (w556, x0, x1_c, x2, x3_c, x4, x5_c, x6_c, x7_c, x9, x10, x11, x13_c, x15, x16, x17_c, x18, x19, x21, x22, x23, x24, x25_c, x26_c, x27, x30, x31_c, x33, x34_c, x36_c, x37, x38, x39_c, x40_c, x42, x43, x44, x45_c, x46, x47_c, x48, x49_c, x51_c, x52_c, x53, x54_c, x55, x56_c, x57_c, x59_c, x60_c, x61, x62, x63, x64, x65, x66, x68_c, x69, x71, x72_c, x73_c, x74_c, x76_c, x77_c, x79, x80, x81, x82, x86_c, x88_c, x89_c, x90, x91_c, x92, x93_c, x96_c, x98_c, x99_c);
and (w557, x0, x2_c, x4_c, x5_c, x7_c, x9, x11, x13_c, x14_c, x15_c, x17_c, x19, x22, x23, x28_c, x32, x33, x36_c, x37_c, x39, x48_c, x50_c, x53_c, x54, x55, x58_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x67_c, x68, x70_c, x71_c, x78, x79_c, x81, x82_c, x83, x85, x86, x87, x89, x90_c, x91_c, x94_c, x95_c, x97, x98_c, x99);
assign w558 = x2_c;
and (w559, x1_c, x3, x4_c, x5, x6_c, x7, x8, x9_c, x11_c, x14, x15, x16, x17, x18, x19_c, x20_c, x22_c, x23_c, x24, x25_c, x27, x28, x29, x30, x31_c, x34_c, x35_c, x36_c, x37, x38_c, x39, x40_c, x41_c, x42, x43, x44, x46_c, x47, x49_c, x50, x51, x52_c, x53_c, x54_c, x55_c, x56_c, x58_c, x59, x60, x63, x64_c, x65_c, x66_c, x68_c, x69, x70, x71_c, x72_c, x73, x78, x79, x80_c, x81_c, x82_c, x83_c, x84_c, x85, x86, x88_c, x89, x92_c, x93_c, x94_c, x95_c, x96_c, x98_c, x99);
and (w560, x0, x1, x2_c, x3_c, x5_c, x9_c, x11, x16, x19_c, x21, x25, x26_c, x27, x28, x30, x32, x33, x34_c, x35_c, x36_c, x37_c, x39, x41_c, x44, x45, x46_c, x50, x51_c, x52, x54_c, x55_c, x56_c, x57_c, x58_c, x60_c, x61_c, x63_c, x64, x66, x67_c, x70, x71_c, x75_c, x79_c, x80, x81, x82_c, x84_c, x88_c, x90, x91_c, x92, x94, x96, x98_c);
and (w561, x3_c, x17, x49_c);
and (w562, x1_c, x10, x15_c, x17, x19_c, x24_c, x27_c, x32_c, x46, x49, x70_c, x75_c, x81, x83_c, x90_c, x98_c);
and (w563, x0, x1, x2, x5, x6, x7_c, x9_c, x10_c, x11_c, x12, x13, x14_c, x16_c, x17_c, x20_c, x21, x24, x25, x26, x27, x29, x31_c, x32_c, x33, x34_c, x37, x38, x40, x41_c, x42_c, x43, x44_c, x46_c, x48, x49, x50, x51_c, x53, x54, x55_c, x57_c, x58, x60, x61_c, x62_c, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x74_c, x75, x76, x77_c, x78_c, x79, x80_c, x81, x82_c, x86_c, x87_c, x88, x89, x90, x91_c, x92, x93, x94, x95, x97_c, x98);
and (w564, x0_c, x1_c, x2_c, x3_c, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14, x15, x17, x18_c, x19, x20_c, x21_c, x22, x23, x24, x25, x26_c, x27_c, x28_c, x29_c, x30_c, x31, x32, x33_c, x34_c, x35, x36, x37, x38, x39_c, x40_c, x41_c, x42, x43, x44_c, x45_c, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55, x56_c, x58_c, x59, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69, x70_c, x71, x72_c, x73, x74, x75, x76_c, x77_c, x78, x79_c, x80_c, x81, x82, x83_c, x84, x85, x86, x87, x89, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97, x98_c, x99);
and (w565, x10_c, x21, x34_c, x44, x45_c, x52, x68_c, x69, x73, x78, x82_c, x83, x88, x94, x99);
and (w566, x2, x4_c, x6, x7, x8_c, x9, x11, x12, x13, x14, x15, x16, x17, x19_c, x20, x21_c, x23_c, x24, x25, x26, x27_c, x28, x29, x31_c, x32_c, x35_c, x36_c, x38_c, x41_c, x42_c, x44, x45, x46_c, x47_c, x50_c, x51, x52_c, x53, x54, x55_c, x56_c, x59, x61, x62, x65_c, x66, x67_c, x68, x69, x71_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x81_c, x82, x83, x84, x85_c, x86, x87_c, x88, x90, x92_c, x93_c, x95_c, x97_c, x98_c);
assign w567 = x73;
and (w568, x0_c, x1_c, x3_c, x4_c, x5, x6_c, x8_c, x9_c, x10_c, x11_c, x13, x14, x15, x16, x17_c, x19, x20_c, x21, x22_c, x23, x24_c, x25_c, x26_c, x28_c, x29, x30, x31_c, x32_c, x33_c, x34, x35_c, x36, x37_c, x39, x40_c, x41_c, x42_c, x43, x44, x46, x47, x48, x50, x51_c, x52, x53, x54_c, x55, x56_c, x57_c, x58_c, x59_c, x61, x62_c, x63_c, x64, x65_c, x66_c, x67_c, x71_c, x72, x73_c, x75_c, x77, x78_c, x79, x80_c, x81, x82, x83, x84, x86, x87_c, x89, x90_c, x92, x93_c, x94_c, x95, x97_c, x98, x99_c);
and (w569, x4, x42_c, x63_c);
and (w570, x0_c, x1_c, x4, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x18, x19, x20_c, x21, x23_c, x26_c, x27, x30_c, x31, x32_c, x33, x34, x35, x38, x42, x48, x49_c, x50_c, x51_c, x53, x56_c, x61_c, x62_c, x66, x67, x68_c, x69_c, x72, x75_c, x76_c, x77_c, x79_c, x80, x81_c, x83_c, x84, x85_c, x86_c, x87, x89_c, x91_c, x93, x94, x95, x96, x98);
and (w571, x0, x3_c, x4_c, x5_c, x6, x7_c, x8_c, x11, x12_c, x13_c, x17, x20, x21, x22, x23, x24_c, x25_c, x27_c, x28_c, x29_c, x30, x31, x32_c, x35_c, x41, x42, x43_c, x45_c, x46, x47_c, x48, x52, x54_c, x55_c, x56_c, x58, x59, x62_c, x63, x64_c, x65, x66_c, x67, x69_c, x70, x71_c, x72, x76, x77_c, x78_c, x79_c, x80_c, x84, x87_c, x91_c, x92_c, x93_c, x95, x96_c, x98_c, x99);
and (w572, x0_c, x2_c, x21_c, x34_c, x38, x60, x78, x83, x84, x86_c, x87);
and (w573, x0, x2_c, x3_c, x4_c, x5, x6, x7, x8_c, x9_c, x10_c, x11, x12_c, x15, x16, x17, x18_c, x19, x20_c, x21, x22_c, x23, x25, x26_c, x27_c, x28, x29, x30, x31, x32, x33_c, x34_c, x35, x36_c, x37, x39, x40_c, x42, x43_c, x44_c, x45, x47_c, x48_c, x49, x50_c, x52, x53_c, x54_c, x55_c, x56, x57_c, x58, x59_c, x60_c, x61, x62_c, x63_c, x64, x66, x67, x68_c, x69_c, x70_c, x71_c, x73_c, x74, x75_c, x78, x79, x80, x82, x85_c, x86_c, x87, x89_c, x90, x91_c, x93, x94, x95, x96_c, x97_c, x98, x99_c);
and (w574, x0_c, x2, x3, x5_c, x6_c, x7, x9, x10, x11_c, x12_c, x13_c, x14_c, x17, x18_c, x20_c, x23_c, x25, x26, x27_c, x29, x30, x31_c, x36_c, x37, x38_c, x39, x40, x41_c, x42, x43_c, x44_c, x46, x47, x48, x49, x50_c, x51, x52_c, x53_c, x54_c, x56, x57_c, x58_c, x60, x61, x62, x63_c, x64, x65_c, x66, x67, x70_c, x72, x74, x75_c, x77, x78_c, x79_c, x81, x82_c, x84_c, x85_c, x86_c, x87, x88_c, x89_c, x90, x91_c, x92, x96, x97_c, x99);
and (w575, x0, x50_c, x51, x53, x67_c, x79, x81);
and (w576, x2, x4, x8_c, x9, x10, x11_c, x12_c, x13, x14_c, x15_c, x16_c, x18, x20, x21_c, x24_c, x25, x29_c, x37, x40, x41_c, x42_c, x43_c, x44_c, x46_c, x49_c, x50, x52_c, x53_c, x55, x56, x58_c, x61_c, x63, x65, x68, x69, x70, x71_c, x73, x74, x76, x77, x78_c, x79, x81_c, x82_c, x83_c, x85, x86_c, x87, x89_c, x91_c, x92, x94_c, x98, x99);
and (w577, x0_c, x1, x2, x3, x4_c, x5_c, x6, x7_c, x8_c, x9_c, x11, x12, x14_c, x15, x16_c, x17, x18, x20_c, x21_c, x22, x23, x25_c, x27_c, x28, x29_c, x30_c, x31, x32, x33_c, x34_c, x35_c, x36_c, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46, x47, x48, x49_c, x50, x51, x52_c, x53_c, x54_c, x55, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x64_c, x67_c, x68, x69, x70, x71_c, x72, x73, x74_c, x75_c, x76, x79, x81_c, x82_c, x83_c, x84_c, x85, x86, x87_c, x88_c, x89, x90, x91_c, x93_c, x94, x95_c, x96_c, x97, x98_c);
and (w578, x0_c, x2_c, x7_c, x12_c, x24_c, x25, x27, x29_c, x30_c, x31, x35, x38, x40_c, x49, x59, x60, x71_c, x72_c, x73_c, x94, x95);
and (w579, x1_c, x2, x5_c, x7, x15_c, x17_c, x18_c, x20, x22_c, x26, x28, x36_c, x43_c, x49, x52, x55_c, x58, x59, x61, x68, x73, x75_c, x77_c, x80_c, x82, x91, x94_c, x95, x96, x98);
and (w580, x0_c, x1, x3_c, x6_c, x7, x8, x10, x12, x13_c, x14, x15, x16, x18, x20_c, x21, x23_c, x24_c, x25, x26, x29_c, x35_c, x37, x39, x41_c, x42_c, x43_c, x44, x45, x48_c, x49, x50, x51, x52_c, x54_c, x55, x56, x57, x59, x61, x62_c, x64, x65, x66, x68_c, x70, x71, x72_c, x75_c, x77, x78, x79, x80, x81, x85_c, x87, x88, x89, x90_c, x91, x93_c, x96, x98_c, x99);
and (w581, x0, x7, x9_c, x12, x13_c, x16_c, x20, x23, x35, x57_c, x58, x70, x75_c, x95);
and (w582, x1, x2, x5_c, x7, x9_c, x12, x13_c, x15_c, x23_c, x26, x28, x30, x38, x40, x45_c, x52_c, x53_c, x55, x59_c, x67, x68, x69_c, x73, x74, x80, x83, x84_c, x89, x90, x92_c);
and (w583, x6, x7, x10, x17, x20_c, x22, x33_c, x45, x46, x50_c, x54, x62, x64, x66_c, x68_c, x71, x73, x74_c, x77, x79, x84, x86_c, x90, x96, x97_c, x99);
and (w584, x0, x1_c, x2_c, x4_c, x6, x9_c, x11_c, x13_c, x14_c, x16_c, x21_c, x23, x24_c, x27_c, x29, x32, x33_c, x36, x37_c, x38_c, x39, x40, x41, x42, x44_c, x45_c, x46_c, x47, x48_c, x51_c, x52, x54, x55_c, x56_c, x58, x61, x62_c, x63, x65_c, x66, x67, x69_c, x70_c, x72_c, x74_c, x75, x77_c, x79, x80_c, x81, x82, x83_c, x84_c, x87, x88, x90, x91, x93, x94_c, x95, x97_c, x98);
and (w585, x2_c, x3, x4, x5_c, x6_c, x7, x9, x12, x13_c, x14, x15, x16, x17, x18, x19_c, x21, x23_c, x25_c, x26_c, x27, x28, x29, x30_c, x32, x33, x34, x35, x36_c, x37_c, x38, x39, x40, x41, x42, x43_c, x44_c, x45, x46_c, x47, x48_c, x49, x50_c, x51_c, x52_c, x53_c, x54, x56, x57_c, x59_c, x60, x61, x62_c, x63_c, x64_c, x65, x66_c, x68_c, x69, x70, x71, x72, x74_c, x75, x76, x77, x78_c, x79, x80, x81_c, x83, x85, x86_c, x87_c, x88, x89_c, x90, x91, x94, x96_c, x97, x98_c, x99);
and (w586, x1_c, x2_c, x4_c, x7, x19, x22, x23, x28_c, x30_c, x33_c, x38, x43_c, x44_c, x52, x64, x72, x74, x76, x79_c, x82, x89_c, x94_c, x95, x99_c);
and (w587, x1_c, x2, x3, x4, x5_c, x6_c, x8, x12_c, x13, x14_c, x15, x16, x17, x18, x20, x21, x23, x27, x29, x30_c, x31, x34, x36, x37, x41_c, x42_c, x44_c, x45, x46_c, x48, x49, x50_c, x51_c, x53_c, x55, x56, x59_c, x61_c, x62_c, x63, x64, x65, x66_c, x69_c, x73_c, x74_c, x75, x76, x77, x80_c, x82_c, x83, x85_c, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x94_c, x97, x98);
and (w588, x0, x1, x2_c, x4, x6_c, x7, x8_c, x9, x10_c, x11_c, x14, x15, x16_c, x17, x18_c, x19, x20, x21_c, x22_c, x23, x24, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31_c, x32, x34_c, x35, x38, x39, x40_c, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48_c, x49, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59, x61_c, x63_c, x65_c, x67_c, x68_c, x69, x70, x72_c, x73, x75, x76, x77_c, x78_c, x79_c, x81_c, x82, x84, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99);
and (w589, x0, x1_c, x2, x3, x4_c, x6_c, x7, x8, x10, x11, x12, x13, x14, x15, x16_c, x17, x19_c, x20, x21_c, x22, x23_c, x24, x25, x27, x28_c, x29, x30_c, x31_c, x32, x33_c, x34_c, x35_c, x36, x37, x38_c, x39, x40, x41_c, x42, x43_c, x44, x46_c, x47, x48_c, x49_c, x50, x51, x52_c, x53, x54_c, x55_c, x57, x58_c, x59, x60, x61_c, x62, x63, x64_c, x65, x66, x67_c, x68, x69, x70, x71, x72, x73, x74_c, x76_c, x77, x78_c, x79_c, x80, x81, x82_c, x83, x84, x85_c, x87_c, x88, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x98, x99_c);
and (w590, x1, x3_c, x6_c, x19_c, x26, x27, x29, x30, x33_c, x39_c, x40, x41, x45_c, x47_c, x52, x58_c, x62_c, x67, x70, x72, x74, x87_c, x88_c, x91_c, x94, x95_c, x97_c, x98_c);
and (w591, x2, x6, x7_c, x9_c, x10_c, x11, x14, x18, x22_c, x23, x24_c, x28_c, x29, x30, x31, x34_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x41_c, x43_c, x44_c, x47_c, x48, x49, x50_c, x51, x53, x55_c, x56_c, x58_c, x59, x62, x63_c, x64_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x75, x77_c, x80, x81_c, x82_c, x83_c, x84_c, x85, x87, x89_c, x90, x91, x93, x96, x97_c, x98_c);
and (w592, x0, x5_c, x6_c, x8, x9_c, x11_c, x12_c, x13, x21_c, x22, x24, x26_c, x28_c, x30, x35, x37_c, x40_c, x41_c, x42, x47_c, x48, x50, x51_c, x53, x55, x56_c, x60, x63, x64_c, x69_c, x80_c, x83, x84_c, x86_c, x88_c, x97_c);
and (w593, x1, x2, x3, x4_c, x5, x7_c, x9_c, x10_c, x11_c, x12_c, x14_c, x16_c, x17_c, x18_c, x19, x20, x21_c, x22, x24_c, x25, x30, x31_c, x32, x37_c, x38_c, x40, x41_c, x42_c, x43, x44_c, x45, x48, x49_c, x50, x52, x53_c, x55, x57_c, x58_c, x59, x61, x65, x69_c, x70, x71, x72_c, x73, x74_c, x75_c, x76, x77, x78, x79_c, x81_c, x82, x86, x87, x88_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c);
and (w594, x27_c, x33, x88_c);
and (w595, x0_c, x1_c, x2, x4, x5, x6, x7_c, x9_c, x10_c, x11, x12, x13, x14_c, x15_c, x16, x17_c, x18_c, x19_c, x20_c, x21, x22, x23_c, x24, x25_c, x27_c, x28, x29_c, x30, x32_c, x33, x37_c, x39, x40_c, x41_c, x43_c, x45_c, x47_c, x48_c, x49, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59, x60, x61, x62_c, x63, x64_c, x65_c, x66_c, x68_c, x69_c, x70, x71, x73, x74_c, x77_c, x78_c, x80, x81_c, x82, x83, x84, x85_c, x86, x88, x90_c, x91_c, x95, x96, x97, x98_c);
and (w596, x1_c, x9_c, x11_c, x15_c, x28_c, x47, x48_c, x49_c, x56_c, x59, x62, x64_c, x75, x78);
and (w597, x2_c, x4_c, x5, x9, x10, x11, x13, x15, x16, x20, x21, x22_c, x23_c, x25, x26_c, x27, x28_c, x31_c, x33, x36_c, x40, x44_c, x47, x52_c, x62, x63, x65_c, x68, x69, x72_c, x73, x74, x76, x78, x81, x83, x84, x85, x87_c, x88, x89, x94, x95);
and (w598, x19_c, x23, x29_c, x37, x40, x44_c, x45_c, x51_c, x65, x67, x73, x95_c, x97_c);
and (w599, x0_c, x3, x4, x7_c, x8, x11_c, x12_c, x14, x30_c, x38_c, x40, x42, x49_c, x50_c, x52_c, x60_c, x73, x74, x75, x77_c, x83_c, x84, x89_c, x90, x97, x98);
and (w600, x0, x1_c, x4_c, x5_c, x6_c, x7_c, x8, x9_c, x10, x11, x13, x15, x16_c, x17, x19, x20_c, x21, x22, x23, x24, x25, x27_c, x28, x29, x30, x31_c, x33, x34, x35, x36_c, x39, x41_c, x43, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50_c, x51, x52_c, x53, x55, x56, x57, x58, x60, x61_c, x63, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x72, x73_c, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81, x82, x83, x84, x85_c, x86_c, x89_c, x91_c, x92_c, x93, x94_c, x95, x96_c);
and (w601, x12_c, x27, x63, x70, x80_c, x88_c, x89, x93);
and (w602, x10, x15, x16_c, x32, x43_c, x52_c, x54, x55_c, x59_c, x63, x71, x81_c, x85_c);
assign w603 = x87_c;
and (w604, x0_c, x2_c, x4_c, x5, x7_c, x11_c, x12, x16_c, x17, x18, x19_c, x24, x25, x33_c, x35_c, x38, x40_c, x41_c, x42_c, x46_c, x47, x48, x50, x51, x56, x57_c, x65, x67_c, x68, x76_c, x81, x87_c, x88_c, x89, x95);
and (w605, x0, x1, x2, x3, x4, x5, x7_c, x8, x9_c, x11, x13_c, x15, x16_c, x18, x19_c, x20_c, x24_c, x25, x26_c, x27_c, x29_c, x30, x31_c, x33_c, x34, x35, x36_c, x37, x38, x39, x41, x43, x45, x47_c, x48_c, x53_c, x55, x57, x58_c, x59_c, x61, x62, x64_c, x65_c, x66_c, x69, x71, x72_c, x74_c, x76_c, x77, x78_c, x81_c, x82_c, x83_c, x84_c, x85_c, x87_c, x88, x89_c, x91, x95_c, x96, x97_c, x99_c);
and (w606, x0, x3, x4, x5, x8_c, x10_c, x12, x13_c, x21_c, x22, x23_c, x25, x26_c, x27_c, x28_c, x29, x33, x36_c, x37, x38_c, x39, x41_c, x42_c, x43, x44_c, x47, x49, x52_c, x55, x57_c, x58_c, x59_c, x61_c, x63_c, x64_c, x66_c, x67_c, x69, x70_c, x71, x72_c, x73_c, x80, x81, x86_c, x90_c, x91, x92, x93_c, x94_c, x95, x97_c, x98);
and (w607, x0, x6_c, x7, x10_c, x11, x12, x13, x15, x18, x19_c, x22_c, x25_c, x26_c, x27, x28_c, x30, x31_c, x33, x34_c, x38, x42_c, x43, x44_c, x46_c, x47_c, x53, x54_c, x55, x56, x57_c, x58, x62_c, x64, x66, x67, x68, x69, x70, x72, x73_c, x74, x75, x81, x83, x85, x89_c, x90, x91_c, x92_c, x96, x98, x99_c);
and (w608, x28, x34, x37, x38_c, x40_c, x44, x46_c, x47, x53_c, x67_c, x69, x73, x76_c, x78, x80_c, x81, x91, x94, x99);
and (w609, x4, x5_c, x9_c, x14_c, x15, x18, x19, x20, x21_c, x23_c, x25, x27_c, x30_c, x32, x33_c, x36, x38, x41_c, x46, x47, x48, x49_c, x50_c, x51, x52_c, x53_c, x59, x61_c, x64, x67_c, x69, x71, x75, x78_c, x81, x83_c, x85_c, x87_c, x89_c, x95);
and (w610, x7, x14, x16, x20, x23_c, x35_c, x42_c, x43_c, x45, x58, x60_c, x64, x65, x69, x82, x85_c, x93_c, x96_c);
and (w611, x1_c, x3, x10, x12, x16, x26_c, x29, x30, x42, x44, x47, x53_c, x54, x57_c, x59_c, x61_c, x68, x69, x74, x81_c, x87, x91);
and (w612, x13, x22, x36_c, x38, x42_c, x54_c, x60, x77, x84, x88_c, x89_c);
and (w613, x0_c, x1, x2, x3, x4, x5_c, x6_c, x7, x8, x9, x10_c, x11, x12_c, x13_c, x15_c, x16, x17_c, x18, x19, x20_c, x21_c, x22_c, x23, x24, x25_c, x27, x28_c, x29, x30, x31, x32_c, x33, x35, x36_c, x37, x38_c, x39_c, x41, x42, x43, x44, x45, x46, x48, x49, x50_c, x51, x52, x53, x54, x55_c, x56, x57_c, x58, x59_c, x61_c, x62, x64_c, x65_c, x66_c, x67_c, x68, x70_c, x71, x72, x74, x75_c, x77_c, x78, x79_c, x81, x82, x83_c, x84, x85, x86, x87_c, x88, x91_c, x92_c, x93_c, x95, x96, x97_c, x98, x99);
and (w614, x0_c, x2, x3_c, x5_c, x6, x7, x10_c, x14_c, x15_c, x17, x20_c, x21, x22_c, x23_c, x24_c, x27, x28_c, x29, x30_c, x31, x34, x36_c, x37_c, x38, x39_c, x41_c, x43_c, x44_c, x46_c, x50_c, x51, x52, x54, x55_c, x57_c, x58_c, x59, x62_c, x63, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x72_c, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x82, x83, x84, x86_c, x87, x88, x89_c, x90_c, x91_c, x92, x94_c, x95_c, x96, x99_c);
and (w615, x0, x5_c, x7, x13, x14_c, x15, x16_c, x19_c, x23, x24, x25_c, x27, x28, x29, x36, x37_c, x39_c, x40_c, x41, x43, x50_c, x51, x55_c, x57_c, x63_c, x64_c, x67_c, x69_c, x73_c, x74, x76_c, x82_c, x90, x91_c, x95, x96);
and (w616, x28_c, x30, x87, x99_c);
and (w617, x21_c, x26_c, x29, x32_c, x56_c, x79_c, x89_c, x94, x95_c, x97, x98_c);
and (w618, x23_c, x71_c);
and (w619, x4_c, x6, x7, x8, x9, x11, x13_c, x14_c, x15, x16_c, x18_c, x20, x21_c, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31, x32, x33, x34_c, x35, x36_c, x37, x39, x40, x41, x42_c, x43, x47_c, x48, x49, x50_c, x52, x53_c, x54_c, x55, x56, x58, x59_c, x61_c, x63, x65_c, x67, x68_c, x69_c, x70, x71, x72_c, x74, x75, x76_c, x77_c, x79_c, x80, x82_c, x83_c, x84_c, x86_c, x90, x91, x93_c, x95, x98);
and (w620, x27, x28_c, x29_c, x34, x45_c, x46, x48, x52_c, x62_c, x82_c, x95, x99_c);
and (w621, x0_c, x5_c, x15, x18, x19, x22, x31, x36, x39_c, x41, x47_c, x49_c, x51, x61, x64, x67, x77, x80_c, x88, x91_c, x96);
and (w622, x0, x1_c, x2, x3, x4_c, x6_c, x7, x8_c, x9, x10, x11_c, x12, x13, x14_c, x15_c, x16_c, x17, x18, x19, x21, x22, x23_c, x24_c, x25_c, x26_c, x27, x29_c, x30, x31, x33, x34, x35, x37, x38, x40, x41, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x53, x54_c, x55_c, x56_c, x59_c, x61, x63, x64, x65, x67_c, x68, x69, x72_c, x73, x74, x75_c, x76_c, x78, x79, x80, x81, x82, x83, x85, x86_c, x87, x88, x89_c, x90, x91, x92, x93_c, x94_c, x95, x96_c, x97, x98_c, x99);
and (w623, x0_c, x1, x2, x6, x7_c, x8_c, x9, x10, x11_c, x12, x14_c, x15, x16_c, x18, x20, x22_c, x23_c, x24_c, x25_c, x26, x27, x31_c, x33, x34, x35, x36, x38_c, x40_c, x41_c, x42, x43_c, x44, x45_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x55, x57_c, x58, x59, x60_c, x61_c, x62, x64, x65, x66, x67, x68_c, x70_c, x73, x74, x75, x76_c, x77, x78, x80, x81, x82_c, x83_c, x84_c, x86_c, x87_c, x89, x90_c, x91_c, x92_c, x94, x95_c, x96, x97_c, x99_c);
and (w624, x5_c, x6, x10_c, x11_c, x19_c, x20_c, x21, x23, x24, x29, x32_c, x34_c, x35, x36_c, x37, x38_c, x39_c, x44, x49_c, x53_c, x55_c, x57, x58, x59, x60, x61_c, x64, x67_c, x68_c, x70_c, x72, x74, x79, x80_c, x81_c, x83, x85, x86, x87_c, x90, x92_c, x96, x98, x99);
and (w625, x69_c, x80_c, x87);
and (w626, x1_c, x2_c, x5_c, x6, x7_c, x9_c, x11, x12_c, x16_c, x17_c, x22, x23, x24, x26, x27, x28_c, x31, x32_c, x36, x37, x38_c, x39, x40, x42_c, x44_c, x45_c, x47, x48_c, x49_c, x50, x51, x52_c, x53_c, x54, x56, x57, x59_c, x61, x62, x65, x66, x67_c, x68_c, x70, x71, x74, x77_c, x78_c, x79, x80, x81_c, x83_c, x84, x85, x86_c, x87_c, x89, x90, x91_c, x92_c, x96_c, x99);
and (w627, x0_c, x8_c, x9, x11_c, x13_c, x14, x17, x18, x22_c, x24_c, x27_c, x30_c, x31_c, x32_c, x35_c, x37_c, x38, x54, x56_c, x58_c, x66, x67, x68, x71_c, x74_c, x77, x82_c, x84_c, x86, x87, x91_c, x98);
and (w628, x1_c, x2_c, x3_c, x6_c, x8, x9, x11_c, x12, x14, x15, x18, x20, x21, x23, x26_c, x27, x29, x31_c, x32, x34_c, x36, x39_c, x40_c, x41, x44, x45, x47_c, x48, x49_c, x52, x53_c, x54, x55_c, x57_c, x58_c, x63_c, x66, x68_c, x69_c, x70, x72_c, x74_c, x75, x77, x78, x83_c, x84_c, x86_c, x87, x89, x91, x92, x93_c, x94, x96_c, x98);
and (w629, x1, x3_c, x4_c, x5_c, x6_c, x7, x9, x10_c, x11, x12_c, x13, x15, x17_c, x18_c, x19, x21, x23_c, x24_c, x25_c, x26, x27, x28, x29, x33_c, x34, x35, x36_c, x37_c, x39, x41_c, x42, x43, x44_c, x45, x49, x51, x52_c, x53, x54_c, x55, x57_c, x59_c, x60, x61_c, x63_c, x64_c, x65, x67_c, x69, x70_c, x71, x73, x75_c, x77, x78, x79_c, x80_c, x81, x82_c, x83, x87, x88_c, x89_c, x91_c, x92_c, x93, x94, x95, x96_c, x98, x99);
and (w630, x0_c, x1, x5, x7_c, x8, x9_c, x10, x11, x12, x13, x14_c, x16_c, x17, x19, x21_c, x22_c, x23, x24, x26, x27_c, x28, x30, x31, x32_c, x34, x35, x36, x37, x38, x39_c, x40, x41, x42, x44_c, x46, x47_c, x48, x49, x50_c, x51, x52_c, x53_c, x54_c, x55, x56, x57, x58, x59, x60, x61_c, x62, x63, x64, x65_c, x67, x68, x69, x71_c, x72_c, x74_c, x78_c, x79_c, x80_c, x81, x82_c, x83_c, x84, x85, x86, x87_c, x88, x89_c, x90_c, x91, x92, x95_c, x96_c, x97_c, x99_c);
and (w631, x1_c, x2, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x12, x13, x14, x15_c, x16, x17, x18_c, x20, x21, x22, x23, x25, x26_c, x28, x30, x31_c, x32_c, x34_c, x35_c, x36_c, x37_c, x38_c, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48_c, x49, x51, x52, x53_c, x54_c, x55, x56_c, x59, x61, x62, x63, x65, x66_c, x67_c, x68, x69_c, x70_c, x73, x74_c, x75_c, x76_c, x77, x78_c, x80_c, x81, x82, x83_c, x84, x85, x86_c, x87_c, x88, x89, x91_c, x92_c, x93, x94, x95, x96_c, x97, x98_c, x99);
and (w632, x0, x1_c, x2, x5_c, x7, x8, x9, x10_c, x12, x13_c, x14_c, x15_c, x16_c, x17_c, x18, x20, x22, x23_c, x24, x25, x26, x27, x28_c, x29, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x38, x39, x40, x41_c, x42, x43_c, x45, x46_c, x47_c, x48_c, x50_c, x51_c, x52, x53, x56, x57_c, x58_c, x59_c, x61_c, x62, x64, x65_c, x66, x67_c, x68_c, x69, x70_c, x71, x72, x73_c, x74, x77, x78, x79_c, x80, x81_c, x82, x84_c, x85, x86, x87, x88, x89, x91_c, x92_c, x93, x94, x95, x96_c, x97_c, x99_c);
and (w633, x11, x12, x18, x20, x23_c, x26, x29, x41_c, x63, x65, x70, x71_c);
and (w634, x0_c, x1, x2, x3_c, x4, x5_c, x6, x7, x8, x9, x10, x11, x12, x13_c, x14_c, x15_c, x16, x17_c, x18, x19_c, x20_c, x21_c, x22, x23, x24, x25, x26, x27_c, x28_c, x29, x30, x31, x32_c, x33, x35_c, x36_c, x37, x38, x39_c, x40_c, x41_c, x42_c, x43, x44_c, x46, x47, x48, x49, x50_c, x51, x52_c, x53, x54_c, x55, x56, x57_c, x58, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70_c, x71_c, x72, x73_c, x74, x75, x76_c, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84, x85, x86_c, x87, x88_c, x89, x90_c, x91, x92_c, x93, x94, x95, x96_c, x97, x98);
and (w635, x0, x1_c, x3_c, x4, x7, x8_c, x10, x12_c, x13, x15, x17, x18, x19_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27, x29, x30_c, x32_c, x34_c, x37_c, x38, x40_c, x41, x42_c, x43, x47_c, x50_c, x51, x52, x53, x54, x55_c, x57_c, x58, x59_c, x61, x62, x63, x65, x66, x67, x69_c, x70_c, x71, x72_c, x73, x74_c, x75, x76, x78_c, x79, x81_c, x83, x86_c, x88_c, x89_c, x90_c, x91_c, x97, x98_c);
and (w636, x1, x2, x3, x5_c, x6_c, x9, x12_c, x13, x14_c, x15, x16, x17_c, x18_c, x19, x20, x21, x24, x26, x27, x28, x29, x30_c, x31, x34_c, x35_c, x36_c, x37_c, x43, x45_c, x46, x47, x49, x50_c, x51, x52, x53_c, x56, x58, x61_c, x62, x65_c, x69_c, x70, x71, x72, x74_c, x75, x76, x77, x78, x81_c, x82, x83_c, x88, x90, x91_c, x92_c, x96_c, x97_c, x98, x99_c);
and (w637, x7, x13, x14, x15_c, x35_c, x37_c, x60, x70, x79, x88, x93_c);
and (w638, x0_c, x1_c, x2_c, x3_c, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11, x12_c, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28_c, x29, x30_c, x31, x32, x33, x35_c, x36, x37_c, x38, x39, x41, x42_c, x43_c, x44, x45, x46, x47, x48_c, x49_c, x50, x51, x52_c, x54, x55, x56, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x66, x67, x68, x69_c, x70_c, x71, x72, x74_c, x75, x76_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87, x88_c, x89, x90, x91_c, x92, x93, x94, x97_c, x98_c, x99);
and (w639, x12_c, x40, x82, x90_c);
and (w640, x4, x5, x9, x15, x19_c, x23, x29, x32_c, x33_c, x38, x40_c, x42_c, x50_c, x62_c, x63_c, x69, x70_c, x73, x74, x79_c, x81, x82_c, x86_c, x91_c, x92_c, x97_c);
and (w641, x0_c, x2_c, x4_c, x5_c, x6_c, x7, x8, x12, x13_c, x14, x15, x16_c, x18_c, x19_c, x22, x23, x24_c, x25, x26, x28, x30, x31, x32, x33_c, x34, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x43, x44, x46, x47_c, x50, x51_c, x52, x53_c, x55_c, x56, x57, x58_c, x60, x62, x65, x66, x67, x68, x69_c, x70, x71, x74_c, x75, x76, x77, x78, x79, x81_c, x84_c, x85_c, x86, x88, x89, x91_c, x93, x95, x96_c, x97_c, x99);
and (w642, x0, x1, x2_c, x3, x4, x5_c, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25, x26, x27, x28_c, x29_c, x30, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43, x44, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56, x57_c, x58, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66_c, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w643, x0_c, x1, x4_c, x5_c, x8, x9_c, x10, x11_c, x13_c, x14, x15_c, x16_c, x17, x18, x19_c, x21_c, x22, x24, x25_c, x28_c, x29_c, x31_c, x32_c, x33, x34, x35, x36, x37, x38_c, x39, x40, x41, x43_c, x47_c, x49, x50, x51, x52_c, x54_c, x55_c, x56_c, x57, x58, x61_c, x62, x63, x64_c, x65, x67_c, x70_c, x73, x74_c, x75, x76_c, x77, x78, x79, x81, x83, x84, x86_c, x88, x89_c, x90_c, x92_c, x93, x98_c, x99_c);
and (w644, x4, x6, x8, x11, x15_c, x16_c, x17, x20, x23, x25_c, x26_c, x29_c, x34_c, x36, x38_c, x41, x47_c, x49_c, x53, x55_c, x64, x67_c, x70_c, x75, x78, x85, x88, x90_c, x91, x92, x95_c);
and (w645, x0, x1, x2, x3, x4, x5_c, x6_c, x7, x8, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x23_c, x24, x25_c, x26, x27, x30, x31, x32_c, x33, x34, x36, x38, x39_c, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48_c, x49_c, x50, x51_c, x52, x53, x54, x55, x56, x57, x58, x59, x60_c, x61_c, x62, x63_c, x64_c, x65, x67_c, x68, x69, x70, x71, x72, x73, x74_c, x75_c, x76_c, x77_c, x78, x80, x81, x82, x83_c, x84, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95_c, x96_c, x97_c, x98, x99);
and (w646, x0_c, x1, x2, x3_c, x4_c, x5, x7, x10, x11_c, x13_c, x15, x18_c, x19_c, x21_c, x23_c, x27_c, x28, x29_c, x30_c, x34, x36_c, x37, x38_c, x40_c, x41_c, x42, x45_c, x47, x48, x49_c, x50, x52_c, x54_c, x56_c, x57_c, x58_c, x62, x63, x65_c, x66_c, x67, x68, x71_c, x74, x75, x77_c, x78, x79, x80_c, x81, x82_c, x88_c, x91, x94, x95_c, x96_c, x98_c, x99_c);
and (w647, x2, x14_c, x15_c, x17_c, x21_c, x22, x25_c, x32_c, x37, x46, x47, x49, x55_c, x56, x57, x60, x71, x72, x80, x83, x86, x88_c, x90, x95_c);
and (w648, x0, x1, x2, x4, x9, x10_c, x11_c, x12_c, x14_c, x15_c, x18_c, x19_c, x21, x25_c, x27, x31, x33, x35_c, x36, x37_c, x38_c, x40, x41, x42, x43_c, x49_c, x50, x53_c, x56, x59, x63, x64_c, x65_c, x66_c, x67, x68, x70, x73_c, x74_c, x75_c, x76, x77_c, x78, x80_c, x81_c, x83_c, x84, x88_c, x89, x90_c, x92, x94_c, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w649, x1, x2, x3, x6_c, x7_c, x8_c, x10, x11, x12, x14_c, x15, x19_c, x20, x21_c, x22, x26, x28_c, x29, x30, x31, x35_c, x36_c, x38, x39, x43_c, x45, x47, x48_c, x52_c, x56, x60_c, x61, x64, x66_c, x69_c, x72_c, x73, x75, x76, x77, x79, x80, x81_c, x83, x93, x95_c, x97_c, x99);
and (w650, x0, x4_c, x6_c, x7_c, x8, x11, x14, x17, x18_c, x19_c, x20_c, x21, x22_c, x24, x25_c, x26, x27, x29, x31_c, x32, x33_c, x35, x36, x38, x39_c, x40, x41_c, x42, x46, x47_c, x48_c, x49_c, x50, x53, x54, x55, x56_c, x57, x58, x59, x60_c, x61, x62_c, x63_c, x64_c, x65_c, x66, x68, x70_c, x73, x74, x75, x76_c, x78, x81, x83_c, x85_c, x88_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x98_c, x99_c);
and (w651, x1_c, x16, x32_c, x49, x64, x80);
and (w652, x0, x1, x2, x3_c, x4_c, x5_c, x7, x8, x9, x10_c, x11, x12_c, x13, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x20_c, x21_c, x22, x23_c, x25, x26, x27, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35, x36_c, x37, x39, x40_c, x41_c, x42, x43, x44_c, x46_c, x47, x48, x49, x50, x51, x52_c, x53_c, x54, x55, x56_c, x57_c, x58_c, x59, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70, x71_c, x74_c, x76_c, x77_c, x78, x79_c, x80_c, x81, x82, x83, x84_c, x86, x87_c, x88_c, x89_c, x90, x91_c, x92, x93, x94, x95, x98, x99_c);
and (w653, x0, x1_c, x2, x3_c, x4, x5_c, x6, x8, x9, x11, x12_c, x13_c, x15_c, x16, x17, x19, x20_c, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34_c, x37_c, x38_c, x39_c, x40_c, x41, x42, x43, x44_c, x45_c, x47, x48, x49_c, x50_c, x51_c, x52, x53, x54_c, x55, x56_c, x57, x58, x59, x60, x61_c, x62, x63, x64, x65, x68, x69, x70, x71_c, x72, x73, x75_c, x77, x79_c, x80_c, x81, x82_c, x83_c, x85_c, x86_c, x87_c, x88_c, x89_c, x92, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w654, x9_c, x14_c, x17, x24_c, x26_c, x56, x61, x73, x79);
and (w655, x0_c, x3, x5, x7, x9, x11_c, x12, x13, x14_c, x16_c, x18_c, x19, x20, x21_c, x22_c, x24_c, x25, x26, x28, x32_c, x34, x35_c, x39_c, x40, x44, x45_c, x46, x47, x48, x49, x50, x51_c, x54, x57, x58_c, x62, x64_c, x65_c, x68, x70_c, x73_c, x76, x77_c, x79, x83_c, x84_c, x85, x87, x89_c, x91, x92_c, x93, x94_c, x96, x97_c, x98, x99_c);
and (w656, x14, x94);
and (w657, x1_c, x3_c, x4, x6_c, x13_c, x21_c, x23, x24_c, x33, x37, x46, x49_c, x54, x55, x57, x58_c, x59, x61, x63, x68_c, x80, x81_c, x89_c, x91_c, x95);
and (w658, x0_c, x4, x7, x8_c, x10_c, x11, x12, x13_c, x14, x15_c, x16, x18, x19, x21_c, x22_c, x25, x26, x27, x29, x30, x31_c, x32, x33_c, x34_c, x35, x37, x46, x48_c, x50_c, x51_c, x52, x53_c, x55_c, x56, x60, x62, x63, x64_c, x65, x66, x67_c, x68, x71, x72, x73, x74_c, x75, x76, x80, x85_c, x88_c, x92_c, x98_c);
and (w659, x1, x2_c, x3_c, x4, x6_c, x9, x10_c, x11_c, x13, x14_c, x16_c, x17_c, x22_c, x24_c, x25_c, x27, x28_c, x29, x30_c, x32_c, x35, x38, x39_c, x43_c, x44, x45_c, x47_c, x48, x49_c, x50, x51_c, x52, x53_c, x56_c, x57, x58, x59, x60, x63_c, x65_c, x66_c, x67, x70, x72, x74, x75_c, x78_c, x79, x80, x81_c, x83, x84_c, x85, x88_c, x89, x90_c, x91, x94, x95_c, x97_c, x99_c);
and (w660, x0_c, x1, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17, x18, x19_c, x20, x21, x22, x23, x24, x25, x26_c, x27_c, x29_c, x30, x31_c, x32_c, x33, x34, x35, x36_c, x37_c, x38_c, x39, x40_c, x41_c, x42, x43, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51, x52, x53, x54_c, x55, x56, x57, x58_c, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69_c, x70_c, x71_c, x72_c, x73_c, x74, x75_c, x76, x77, x78, x79, x80, x81, x82, x83_c, x84_c, x85_c, x86, x87, x88_c, x89_c, x90, x91, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w661, x1_c, x2, x4, x6_c, x7, x8, x10, x12, x18, x20, x21, x22_c, x23_c, x24, x25_c, x26_c, x27_c, x30, x31_c, x32_c, x36_c, x39, x42_c, x44_c, x46, x47_c, x48, x49_c, x51_c, x54_c, x55, x56, x57, x58_c, x66, x69_c, x71, x72, x75_c, x79, x82_c, x83, x84_c, x85, x88, x89_c, x90_c, x92_c, x95, x96_c);
and (w662, x4, x5, x6_c, x7, x8_c, x9_c, x10, x12_c, x13_c, x14_c, x15_c, x16, x17, x18, x19, x20_c, x21, x22_c, x23_c, x24, x26_c, x27_c, x28, x29, x30, x31_c, x32, x33_c, x34, x35_c, x36, x38, x39_c, x40, x41_c, x42_c, x43_c, x45, x46, x48_c, x49_c, x50, x52, x53, x54, x55_c, x57, x58, x59_c, x60_c, x61_c, x62, x63_c, x64, x66, x67, x68_c, x69, x71, x74_c, x75_c, x76, x77_c, x78_c, x81_c, x82_c, x83, x84_c, x85_c, x86_c, x87_c, x88, x89, x90_c, x92, x94, x95_c, x96, x97_c, x98_c, x99);
and (w663, x0_c, x16, x38, x53_c, x84, x99);
and (w664, x0, x1_c, x5_c, x6, x7_c, x8, x9, x10, x11, x12, x14, x15_c, x16_c, x17_c, x18_c, x19_c, x20_c, x23, x24_c, x27, x28, x29_c, x30, x32_c, x36, x37_c, x40, x41_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49, x50, x51, x52, x53_c, x54, x55, x56_c, x57_c, x58_c, x59, x62_c, x64, x65, x66, x67, x68, x69, x70, x71_c, x72_c, x73_c, x74, x77, x78, x79, x81_c, x83, x85, x86, x87_c, x88_c, x89, x90_c, x91, x93_c, x94, x95_c, x96_c, x98_c);
and (w665, x87, x96);
and (w666, x0_c, x3, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x11, x12, x15, x16_c, x17, x18_c, x19_c, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x28_c, x29, x30, x31_c, x32, x33, x34_c, x35_c, x36, x37_c, x38, x39, x40, x41_c, x42_c, x43_c, x44, x45_c, x46_c, x48, x49, x50, x51, x52, x53, x54_c, x55, x56, x57_c, x58_c, x59_c, x60, x61_c, x62_c, x63_c, x64, x65, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x73_c, x74, x75, x76, x77, x78_c, x79, x80_c, x81, x82, x83_c, x84, x87, x89_c, x90_c, x91_c, x92, x93, x94, x95, x96, x97_c, x98, x99_c);
and (w667, x4, x5, x7_c, x10_c, x11_c, x18, x19, x21_c, x22, x28, x29, x30, x31_c, x32_c, x35_c, x36, x37_c, x38, x45_c, x49, x51, x52, x53_c, x55, x59, x62_c, x64_c, x67, x69_c, x70, x74_c, x75, x78, x79, x80_c, x81, x83_c, x86_c, x87_c, x90, x94, x95, x96, x97);
and (w668, x2, x5_c, x7, x28_c, x32_c, x33_c, x36, x41_c, x57, x62_c, x73_c, x75, x80_c);
and (w669, x0_c, x1, x2, x3_c, x5, x6, x7_c, x8, x9_c, x10_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28_c, x29_c, x30, x31_c, x32, x34, x35_c, x37, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45, x46_c, x47, x49, x50_c, x51_c, x52_c, x53_c, x54, x56, x58_c, x59_c, x61, x62_c, x63, x64, x65, x66, x67, x68_c, x69, x70_c, x71, x72_c, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84, x85, x86, x87_c, x88, x89, x90, x91, x92_c, x95, x96, x97_c, x98, x99_c);
and (w670, x0, x1_c, x2_c, x4, x5, x6, x8_c, x9_c, x10_c, x13, x14, x15_c, x16_c, x17_c, x19_c, x20, x21_c, x23_c, x24, x25, x32, x34, x35_c, x39, x41, x42, x44_c, x45, x46_c, x47, x49_c, x54_c, x55_c, x56, x57_c, x61, x62_c, x64_c, x68, x70, x71_c, x72_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82_c, x83_c, x85, x86_c, x87, x88, x89_c, x91_c, x92, x93, x94, x95, x96, x97_c, x99);
and (w671, x0_c, x6, x10, x17_c, x29_c, x52, x58_c, x74_c, x89, x92_c, x96, x97);
and (w672, x0, x1_c, x2, x3_c, x4, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12_c, x13, x15, x17_c, x18, x19, x20_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x34, x35, x36, x37_c, x38_c, x39, x40, x41_c, x43, x44_c, x45_c, x46, x47, x48, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x56, x57_c, x58_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x66, x67, x68_c, x69_c, x70, x71, x72, x73_c, x74_c, x75_c, x76, x77, x78, x79_c, x80_c, x81_c, x82, x83, x84, x85_c, x86_c, x87, x88, x89_c, x90, x91, x92_c, x93, x94, x95, x96, x97, x98_c, x99_c);
and (w673, x0_c, x2, x5, x8, x12_c, x14_c, x18_c, x22_c, x24_c, x25_c, x27, x33, x40_c, x47_c, x48, x52, x54_c, x55_c, x61, x62, x63, x70_c, x74_c, x79_c, x80, x84, x85_c, x86_c, x87, x89_c, x91, x92_c, x93_c, x94, x95_c, x96, x99);
and (w674, x21, x30, x39_c, x50_c, x54_c, x64, x71_c);
and (w675, x0, x2_c, x3_c, x5_c, x7_c, x8, x9, x13_c, x16, x17_c, x20, x21, x23, x24, x25_c, x29_c, x32, x33_c, x34_c, x35, x39, x40_c, x41_c, x42, x44_c, x45, x46_c, x48_c, x49, x51_c, x52, x53, x55_c, x56, x58_c, x59_c, x60, x62, x65, x66, x67_c, x70, x71, x72_c, x73, x74, x75_c, x76_c, x77_c, x79, x80_c, x86_c, x89, x93_c, x96, x99);
and (w676, x1, x2_c, x6, x7_c, x8, x9, x10, x11_c, x12_c, x13_c, x14, x16_c, x17_c, x19, x20_c, x21_c, x22, x24_c, x31, x33_c, x35, x36_c, x37_c, x38, x39_c, x40_c, x42, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x58_c, x59_c, x61_c, x62, x63, x64_c, x66_c, x67_c, x69, x71_c, x72_c, x73_c, x74_c, x75, x77, x78, x82, x84_c, x85, x88, x89_c, x90, x91_c, x92_c, x93, x96_c, x97, x98, x99_c);
and (w677, x0, x6_c, x12, x13_c, x15_c, x17_c, x18_c, x19_c, x20, x22_c, x23, x25_c, x29_c, x30, x32, x35, x40_c, x41_c, x45_c, x46, x47, x49_c, x50, x52, x56, x58_c, x60_c, x62, x64, x65, x66, x68, x71_c, x72_c, x76, x77, x78, x79_c, x88_c, x89_c, x90_c, x91, x92, x93_c, x97_c, x99);
and (w678, x1_c, x41, x55, x65_c, x74_c, x89, x94_c);
and (w679, x3_c, x5, x6, x7_c, x10, x12_c, x13, x14_c, x19_c, x20_c, x26_c, x29_c, x30_c, x32, x34_c, x35, x36_c, x42_c, x43, x44, x46, x47, x49, x50, x51_c, x53_c, x54_c, x56, x57, x61_c, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x70_c, x73, x74, x80, x82_c, x83_c, x84, x85, x87_c, x88_c, x89_c, x90, x92_c, x94_c, x95_c, x97_c, x99_c);
and (w680, x0, x2, x4, x5_c, x6, x8, x9_c, x12, x13, x15_c, x16, x17_c, x18_c, x19, x22_c, x23_c, x25_c, x27_c, x28, x29_c, x30_c, x31_c, x33_c, x35_c, x36, x38, x40, x41, x42_c, x43_c, x45_c, x46, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x56_c, x58, x61_c, x62, x63, x65, x68, x69_c, x70, x71_c, x73, x75, x76_c, x78_c, x79_c, x80, x82_c, x83_c, x86_c, x90, x91, x92_c, x93, x94_c, x96, x97);
and (w681, x1_c, x3_c, x5, x7, x9, x11_c, x12_c, x13_c, x15_c, x16, x17, x18_c, x19_c, x20_c, x21, x24_c, x26, x27, x30, x31, x33, x36_c, x37_c, x38_c, x39_c, x40_c, x42, x43_c, x45, x48_c, x51, x52, x56_c, x57_c, x58_c, x60, x61_c, x62, x63_c, x64_c, x66, x67_c, x68, x72, x73, x74, x75_c, x76, x77_c, x78_c, x80_c, x81_c, x83, x85, x86, x87, x90_c, x92, x94, x97, x98_c);
and (w682, x1_c, x2, x3, x6_c, x7, x8, x9_c, x11, x15, x16, x18, x19_c, x21, x22, x23, x25, x27_c, x30_c, x31_c, x32, x35, x36_c, x37_c, x38_c, x39_c, x41, x42, x44, x45_c, x46_c, x47, x48_c, x50, x51, x52, x53_c, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61_c, x62, x63_c, x65, x66, x67_c, x68, x70, x71, x73_c, x74, x75, x76, x77, x78_c, x79_c, x81_c, x82_c, x84_c, x87, x88, x92_c, x93_c, x95_c, x96, x97, x98, x99);
and (w683, x1_c, x3, x4, x5_c, x6_c, x7_c, x8_c, x9, x10, x12_c, x13, x14, x15_c, x16_c, x17, x18, x20_c, x21, x22, x23, x24, x25, x26_c, x28, x30, x32_c, x33_c, x35, x36_c, x39, x40_c, x41, x44_c, x45, x47_c, x48, x49_c, x50, x54_c, x55_c, x57_c, x59, x61, x63, x64, x65_c, x66_c, x67, x69, x71, x73, x74, x75, x77_c, x79, x80, x81_c, x82, x83, x85_c, x88, x89_c, x90, x91_c, x93_c, x96, x97, x98_c, x99_c);
and (w684, x0, x1, x2, x5, x7, x9_c, x11, x12, x13_c, x14, x16, x17, x18, x19, x20, x21, x22_c, x24, x26_c, x29, x30_c, x31_c, x32_c, x33, x34, x36, x37, x38, x40_c, x41_c, x43, x46_c, x47_c, x48, x49, x50, x51, x52, x55_c, x57, x59_c, x60_c, x61, x65_c, x66, x69_c, x70_c, x71_c, x72, x73, x74_c, x78_c, x80, x81_c, x83_c, x84_c, x86, x88, x89, x90, x91_c, x93_c, x94, x95_c, x97_c, x99_c);
and (w685, x3, x5_c, x7_c, x8_c, x11_c, x14_c, x15_c, x16_c, x17, x18_c, x20, x21, x22_c, x24_c, x29_c, x30_c, x31_c, x32, x33, x34_c, x39, x41, x52_c, x54, x55, x56_c, x57_c, x58, x63_c, x64, x68_c, x69_c, x79_c, x82_c, x83_c, x84_c, x86_c, x88, x89, x90_c, x95, x96, x97_c);
and (w686, x1, x2_c, x6_c, x15, x16, x47, x57, x79_c, x95_c, x97);
and (w687, x0_c, x1_c, x2_c, x3, x4, x5, x6_c, x7_c, x8, x9_c, x10, x11, x13, x14, x16, x17_c, x20, x21, x23, x24, x27, x28, x29, x32, x34, x35_c, x36_c, x37, x38_c, x39_c, x42, x43, x46_c, x47, x48_c, x49, x50, x51_c, x52, x53_c, x54, x55, x56_c, x58, x59, x60, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69_c, x70, x72_c, x76, x78_c, x79_c, x80, x82, x83_c, x85_c, x87, x89, x90_c, x91_c, x92_c, x93, x94_c, x95, x96, x98, x99);
and (w688, x0, x1, x2, x3, x4_c, x6_c, x7, x10, x11_c, x13, x14_c, x15, x16, x17_c, x18, x20_c, x21_c, x22_c, x23_c, x25, x26, x27, x29_c, x30_c, x31, x35_c, x36, x37_c, x39, x40, x41, x42, x43_c, x45, x46_c, x47_c, x49_c, x52_c, x54, x58_c, x59, x60, x61, x62, x64_c, x65_c, x68, x69_c, x70_c, x71, x72, x73, x74, x76_c, x77_c, x78_c, x82, x83, x84_c, x86_c, x87_c, x88_c, x89, x90_c, x91, x92, x96_c, x97_c, x98, x99);
and (w689, x0_c, x1_c, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11_c, x12_c, x13, x14, x15_c, x16, x17, x18, x19_c, x20, x21, x22, x23_c, x24_c, x25, x26_c, x27_c, x28, x29, x30_c, x31, x32, x33, x34_c, x35_c, x36_c, x37, x38_c, x39, x40, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52_c, x53, x54, x55_c, x56_c, x57_c, x58_c, x59, x60_c, x61, x62_c, x63, x64, x65, x66, x67, x68, x69, x70, x71_c, x72_c, x73_c, x74, x75_c, x77_c, x78_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90, x91_c, x92, x93_c, x94, x95_c, x96, x97_c, x98_c, x99);
and (w690, x0, x2_c, x5_c, x12, x13, x14_c, x16, x24, x25_c, x26, x30, x33_c, x34_c, x40_c, x43, x44_c, x45, x46, x53_c, x58, x59_c, x61, x63_c, x68, x69, x75_c, x77, x78, x79_c, x80, x81, x83_c, x85, x87, x89, x90, x92, x93_c, x94_c, x98);
and (w691, x38, x39, x84_c);
and (w692, x36_c, x48_c, x63_c, x80_c);
and (w693, x0, x1, x2_c, x4_c, x7_c, x10_c, x13_c, x15_c, x18_c, x20_c, x23_c, x27_c, x28, x29_c, x31, x35, x37, x41, x42, x44_c, x46, x48_c, x49_c, x50, x55_c, x56_c, x57, x58_c, x60_c, x64, x66, x68_c, x73_c, x74, x75_c, x76_c, x78, x79_c, x82, x83, x85_c, x86_c, x90_c, x93, x94, x95_c);
and (w694, x0_c, x1_c, x3_c, x4_c, x5_c, x6, x7_c, x8, x9_c, x11_c, x12_c, x13_c, x15_c, x16, x17_c, x18_c, x20, x23, x24_c, x25, x26, x27_c, x28, x29, x30, x33, x34, x36, x37, x38_c, x43_c, x45_c, x46_c, x47, x49_c, x50, x51, x52_c, x54_c, x55_c, x56_c, x58, x60_c, x61, x62_c, x63_c, x64_c, x65, x66, x67, x68, x69, x70, x71, x73, x74, x79_c, x82, x84, x85, x86, x88_c, x89, x91, x93_c, x94, x96_c, x97, x98_c);
and (w695, x0_c, x2, x5_c, x6, x7_c, x9_c, x10, x13_c, x14_c, x15_c, x16, x17, x18, x20, x21_c, x22_c, x23, x25_c, x26, x27, x28, x29_c, x31_c, x32_c, x33, x35_c, x36, x37_c, x38_c, x39_c, x40, x42_c, x45, x47, x48, x49_c, x51_c, x52, x55, x56, x57, x58_c, x61, x64, x67, x68, x70_c, x71, x72, x73, x74, x75, x77, x78_c, x79_c, x81, x82, x84_c, x85, x86_c, x87, x88_c, x89_c, x91_c, x92_c, x93, x94, x97);
and (w696, x0, x1, x2, x3_c, x4, x6_c, x7_c, x8_c, x9, x10, x11_c, x12, x13, x14_c, x15, x18, x19, x20_c, x22_c, x23_c, x24_c, x25, x26, x28_c, x29, x32_c, x33, x34_c, x35_c, x36, x37, x38, x40, x42, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x51, x52, x53_c, x54_c, x55, x56_c, x57_c, x58, x59, x60_c, x61, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68_c, x71, x72, x74_c, x75_c, x76_c, x77, x79_c, x81, x82, x83_c, x84, x85, x86, x87, x88, x91, x92_c, x93, x96_c, x97_c, x98_c, x99);
and (w697, x22, x34_c, x55, x63_c, x76_c, x80, x91);
and (w698, x12_c, x32, x91);
and (w699, x12_c, x29, x46, x47_c, x48_c, x50_c, x61_c, x66, x67_c, x77, x78, x94);
and (w700, x2_c, x3_c, x5, x7, x8, x9_c, x10_c, x12, x13, x16, x17, x20_c, x22_c, x24_c, x26_c, x27_c, x28, x29_c, x30_c, x31_c, x32, x33_c, x35_c, x36, x41_c, x42, x43, x44, x45_c, x46, x47, x50, x51, x52, x53, x57_c, x58_c, x60_c, x62_c, x63, x64, x65, x66, x69_c, x72_c, x73, x76, x78, x80, x81_c, x83, x85_c, x87, x89_c, x95, x98_c, x99_c);
and (w701, x0, x2, x3, x6_c, x10_c, x11, x13_c, x21, x24, x25, x33, x38_c, x44_c, x57, x65_c, x67_c, x69, x72_c, x74_c, x77_c, x81, x91, x98_c);
and (w702, x0, x1, x3, x5_c, x7_c, x8_c, x10_c, x11, x12_c, x13, x17, x18_c, x19, x21_c, x22, x23, x25, x30_c, x34_c, x35_c, x36_c, x37_c, x39_c, x42_c, x43, x44_c, x45, x46_c, x49_c, x51_c, x52_c, x53, x57, x59, x60_c, x61_c, x64_c, x68, x69, x70_c, x72_c, x73, x74_c, x75, x76_c, x79, x81, x84_c, x88, x89_c, x92_c, x93_c, x96);
and (w703, x0_c, x1, x2, x3_c, x4, x5, x6, x7, x8_c, x9, x10_c, x11, x12, x13, x14, x16_c, x18_c, x19_c, x20, x21_c, x22_c, x23, x24_c, x25, x26_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34, x36_c, x37, x38, x40, x41_c, x42, x44_c, x45_c, x46_c, x47_c, x48, x49_c, x50, x51_c, x54_c, x55, x56_c, x58_c, x60_c, x61_c, x63_c, x65_c, x66, x68, x70_c, x71, x72, x74_c, x76_c, x77, x79, x81_c, x82_c, x83, x84, x85, x86_c, x88_c, x90, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98_c, x99_c);
and (w704, x0, x6_c, x7_c, x9, x12_c, x14, x15, x17, x19, x20_c, x22_c, x23_c, x25, x26, x27, x28_c, x30_c, x34_c, x36, x37_c, x42, x43, x46, x47, x49_c, x53_c, x55, x56_c, x58_c, x61_c, x62_c, x64, x65_c, x67_c, x69_c, x74_c, x76, x77, x78_c, x81, x82, x83_c, x84_c, x86_c, x87_c, x89_c, x91_c, x92_c, x94, x95, x96_c, x98_c, x99_c);
and (w705, x7_c, x22_c, x28_c, x40, x41_c, x43_c, x45, x54_c, x63);
and (w706, x0, x1_c, x2, x3_c, x4_c, x5, x6, x7, x8, x9, x11_c, x12_c, x13, x14, x15, x16_c, x17, x18, x19_c, x20_c, x21, x22_c, x23_c, x24_c, x25_c, x26, x27_c, x28_c, x29_c, x30, x32, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x40, x41, x42, x44_c, x45_c, x47, x48_c, x49, x50, x51, x52, x53_c, x54, x55, x56_c, x57_c, x58_c, x59_c, x60, x61_c, x62, x63, x64, x66, x67, x68, x69_c, x70_c, x71_c, x72, x73, x74, x75_c, x76_c, x77, x78_c, x79_c, x80, x81_c, x82_c, x83, x84_c, x85, x86, x87, x88_c, x89_c, x90, x91, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w707, x1_c, x3, x8, x11_c, x12, x13_c, x15_c, x16, x18, x20_c, x21_c, x23_c, x25_c, x26, x28, x29_c, x31, x33_c, x37_c, x39_c, x40_c, x43_c, x44, x45_c, x46_c, x48_c, x51, x53, x54, x58_c, x59, x62_c, x63, x64_c, x65, x66_c, x69_c, x72, x75_c, x79_c, x80, x83_c, x84_c, x86_c, x96_c, x97, x98_c);
and (w708, x0, x1_c, x3_c, x5_c, x6, x8, x9, x10_c, x11, x12, x15, x16_c, x17, x18, x19, x20, x21_c, x22, x23_c, x25_c, x27_c, x28_c, x29, x30_c, x31, x32_c, x34, x35, x36_c, x38, x39_c, x40_c, x41_c, x43, x44, x45, x47_c, x48_c, x50_c, x53_c, x55, x56, x58, x60, x61, x62, x64, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x74_c, x76_c, x77, x78_c, x79, x81, x82_c, x84, x85_c, x86, x87, x88, x89_c, x90, x91, x92, x93_c, x94, x95, x97_c, x98_c, x99);
and (w709, x0_c, x1_c, x2_c, x9_c, x10_c, x12, x13, x21_c, x25, x26_c, x27_c, x34_c, x39_c, x45_c, x48, x53, x55, x56_c, x60, x64, x70_c, x72, x74_c, x76_c, x78_c, x79_c, x80, x82_c, x84_c, x85_c, x88, x89, x90, x94_c, x95, x98_c, x99);
and (w710, x0, x1_c, x3_c, x4, x5, x6_c, x7, x8_c, x9_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x18_c, x19, x20_c, x21, x22, x23, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32_c, x33, x34, x35_c, x37, x38, x39, x40_c, x41_c, x42_c, x43_c, x45_c, x46, x47, x48_c, x49_c, x50_c, x51_c, x52_c, x53_c, x54_c, x55_c, x57_c, x58_c, x59, x60, x61, x62_c, x63, x64_c, x65, x66_c, x68_c, x69, x70_c, x71, x72, x73, x74_c, x75, x76, x77_c, x78_c, x79, x80, x81_c, x83_c, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99_c);
and (w711, x0, x1_c, x2_c, x3, x4_c, x5_c, x6, x7, x8, x9, x10_c, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x18, x19, x20, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34_c, x35, x36, x37_c, x38_c, x39, x40_c, x41, x42_c, x43, x44, x45, x46_c, x47_c, x48, x49, x50, x51_c, x52_c, x53_c, x54, x55_c, x56_c, x57, x58_c, x59, x60, x61_c, x62_c, x63, x64, x65_c, x66_c, x67_c, x68_c, x69, x70, x71_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78_c, x79_c, x80, x81, x82, x83, x84_c, x85_c, x86_c, x87, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w712, x1_c, x2, x4, x5, x6_c, x8_c, x9, x11_c, x13, x14_c, x16_c, x19, x20_c, x21, x22_c, x23_c, x24, x25, x26_c, x27_c, x29_c, x30_c, x31, x33, x34_c, x35, x36, x40, x41_c, x42_c, x43, x44, x45, x46, x47, x48, x50_c, x52_c, x53, x55_c, x57_c, x59, x61_c, x62_c, x63_c, x65_c, x66, x67, x70, x71, x72, x73_c, x74, x75, x76_c, x77_c, x79, x82, x83_c, x85_c, x90, x91, x92, x94_c, x95_c, x96, x97_c, x98_c, x99);
and (w713, x0_c, x5, x7, x12_c, x13, x14, x16_c, x19, x20, x24, x27, x29_c, x31, x33_c, x36, x37, x38, x40, x41_c, x42_c, x43, x44_c, x45_c, x47_c, x50_c, x53, x65, x67_c, x68, x69_c, x70, x71, x75, x78_c, x79_c, x81_c, x82, x83_c, x84_c, x86_c, x92, x93_c, x94, x95, x96_c, x98);
and (w714, x1_c, x3_c, x6, x9, x10, x13, x14_c, x17_c, x18, x19, x21_c, x22_c, x23_c, x24_c, x27, x28_c, x29_c, x30, x31_c, x36, x38_c, x39_c, x40_c, x41, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x52, x54, x57_c, x58, x59, x60, x62, x64_c, x67, x68_c, x70_c, x72, x74_c, x75_c, x76_c, x77_c, x78_c, x80_c, x81_c, x82, x84_c, x87_c, x89, x90, x92_c, x93, x94_c, x96_c, x97, x98);
and (w715, x10_c, x11, x13, x15, x17, x20, x27_c, x31_c, x44, x46, x55_c, x68, x78_c, x81, x88_c, x91_c, x93_c);
and (w716, x0, x1_c, x2, x3, x4, x5, x6_c, x7, x8_c, x9_c, x10, x11_c, x13_c, x14, x15_c, x16, x17_c, x19_c, x20_c, x22_c, x23, x24_c, x25, x26_c, x28, x29_c, x30, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37, x38, x39_c, x40, x41_c, x43, x44, x45, x46, x47_c, x48, x49_c, x50_c, x51_c, x52, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61, x62, x63, x64, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x72_c, x73_c, x74_c, x75_c, x76_c, x77, x78, x79_c, x80, x81_c, x82, x83, x84, x85_c, x86, x87, x89, x90, x91, x92_c, x93, x94_c, x95, x96, x97_c, x98, x99_c);
and (w717, x2_c, x4_c, x9_c, x11, x15, x16_c, x21, x25, x33_c, x37, x40_c, x45, x47, x54_c, x55_c, x67, x68, x69_c, x71, x81_c, x82, x88_c, x93_c, x95_c);
and (w718, x0_c, x2_c, x3_c, x4, x6, x7, x8, x11_c, x13, x14, x15_c, x16, x17, x18, x21_c, x26_c, x27, x28, x30_c, x31_c, x32, x34, x35, x36_c, x38, x40, x43, x47_c, x48_c, x53, x54, x55_c, x57, x58_c, x63_c, x65_c, x66, x68_c, x69, x70_c, x71, x75, x76, x77, x78_c, x79, x80_c, x83_c, x84_c, x85, x87_c, x90, x92, x93_c, x97_c, x98, x99_c);
and (w719, x0, x3, x4, x8_c, x11_c, x12, x13_c, x14, x17_c, x18_c, x19, x22_c, x23_c, x26_c, x27, x28, x29_c, x30, x31, x33, x34_c, x36_c, x37, x38, x40, x43_c, x45_c, x47_c, x48_c, x49, x50_c, x51_c, x52, x53_c, x57, x58_c, x60, x64, x68, x71_c, x74_c, x75, x78_c, x79_c, x80, x83_c, x84, x86_c, x89_c, x92, x93_c, x94_c, x95_c);
and (w720, x3_c, x4, x5_c, x7, x25_c, x36, x38, x46_c, x49, x51_c, x54, x61, x63_c, x76_c, x77_c, x78, x89, x91, x93);
and (w721, x23, x46_c, x51_c, x58);
and (w722, x1_c, x6_c, x14, x29_c, x49);
and (w723, x2_c, x10, x15, x24_c, x26_c, x27, x28, x35_c, x39, x46, x48, x50, x51_c, x58_c, x61_c, x64_c, x66_c, x69_c, x73_c, x74_c, x76, x81_c, x82, x84, x86_c, x88, x89, x98, x99_c);
and (w724, x8, x18, x20_c, x40, x66, x78, x80_c, x82_c);
and (w725, x9_c, x10_c, x12, x15_c, x16, x25_c, x26_c, x27_c, x34, x36, x37, x39_c, x42_c, x56_c, x59_c, x86_c, x88, x93, x95, x98_c);
and (w726, x0_c, x1, x2_c, x3_c, x5, x6, x9, x11_c, x12_c, x13_c, x14_c, x15_c, x18_c, x19_c, x20, x21_c, x24_c, x25, x26, x29, x30_c, x32, x34_c, x35, x36_c, x37_c, x40, x41, x43_c, x44, x48_c, x50_c, x51, x52_c, x53, x56, x57, x60, x62, x64, x66_c, x67_c, x69, x71_c, x72, x74, x75, x76, x80, x86_c, x88, x89_c, x92_c, x98_c, x99_c);
and (w727, x0, x2_c, x5, x6, x12, x15, x20_c, x24_c, x28, x31, x33_c, x35_c, x36_c, x37, x38_c, x44_c, x46, x47_c, x50, x51_c, x52_c, x55_c, x56, x58_c, x65, x69, x72, x73, x83_c, x90_c, x92, x99);
and (w728, x0, x1, x2_c, x3, x4_c, x5_c, x6, x8_c, x9, x10_c, x11_c, x12_c, x13_c, x15_c, x16_c, x17, x18, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x29_c, x30_c, x34_c, x35, x36, x37, x38, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47, x48_c, x49_c, x50, x51_c, x52_c, x53, x57, x58_c, x59, x60_c, x61_c, x62, x63, x64_c, x65, x67, x68_c, x71_c, x72_c, x73, x74, x75, x77, x78_c, x79_c, x81_c, x82, x84_c, x85_c, x87_c, x88, x89_c, x90, x91, x92, x93_c, x94, x96, x98_c, x99);
and (w729, x2, x3, x4, x5_c, x6, x7, x8_c, x9, x10_c, x11, x12_c, x13_c, x14_c, x15_c, x16_c, x18, x20_c, x21, x22, x23, x24, x25_c, x26_c, x27_c, x28, x29, x32, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x47, x48, x50, x51, x54_c, x55, x56, x57_c, x58, x59, x60_c, x61_c, x62_c, x63_c, x64_c, x65_c, x66_c, x67, x68, x69, x70_c, x72_c, x73_c, x74, x75, x76_c, x77, x79, x80_c, x81, x82, x83, x84_c, x85_c, x87_c, x88, x92, x94_c, x95_c, x96, x97_c);
and (w730, x11_c, x27, x37, x50, x51, x55_c, x57, x59, x64, x66_c, x71, x75_c, x76, x79_c, x86_c, x99_c);
and (w731, x2, x4_c, x7, x9, x10, x13, x14, x15, x16, x17_c, x18_c, x19_c, x20, x24_c, x26, x27, x29, x30, x32_c, x35, x36, x37, x40_c, x41, x43_c, x46_c, x48, x50_c, x52_c, x53_c, x55, x56_c, x60_c, x62, x66_c, x67_c, x69, x73, x75, x76, x77, x78_c, x79, x82, x83, x84_c, x85, x86, x87, x89_c, x91, x92_c, x93_c, x94_c, x97_c, x99);
and (w732, x2_c, x3, x4, x7, x11_c, x13_c, x16, x18_c, x19_c, x21_c, x26, x35, x37, x38_c, x41, x44_c, x52_c, x56, x57, x60_c, x62, x68, x70, x75_c, x76, x82_c, x83, x91, x96, x98);
and (w733, x0, x1, x2, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x12_c, x13_c, x15, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28, x29, x30_c, x31, x32_c, x33_c, x34_c, x35, x36, x38_c, x39, x40_c, x41, x42, x43_c, x44_c, x45, x46, x47_c, x48, x49_c, x50, x51, x52_c, x53_c, x55_c, x56_c, x57_c, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64, x65_c, x66_c, x67_c, x68, x70, x72_c, x73, x74_c, x78, x79, x81, x82_c, x84_c, x86, x87_c, x88, x90, x91_c, x94, x95, x97_c, x98, x99);
and (w734, x6, x26_c, x34_c, x41, x44_c, x49_c, x60, x71, x77_c, x90_c, x93_c);
and (w735, x3, x5_c, x6_c, x7_c, x9, x11_c, x12, x14_c, x15_c, x18, x19_c, x20, x21, x22_c, x25_c, x29_c, x30_c, x38, x39_c, x41, x44_c, x46, x47, x48_c, x50_c, x52_c, x53_c, x55_c, x57, x58, x59, x61_c, x62_c, x63_c, x70, x73_c, x74_c, x78_c, x82, x85_c, x86_c, x87_c, x88, x90, x92, x95, x96_c, x97, x98_c);
and (w736, x1, x2_c, x3, x4_c, x7, x8_c, x9, x13_c, x14_c, x15, x17, x18_c, x24_c, x26, x31_c, x33, x35, x36_c, x38, x39, x40, x41_c, x42_c, x43, x44_c, x50_c, x52, x56_c, x58_c, x62_c, x65_c, x67, x70, x72_c, x73_c, x75, x76_c, x77_c, x79_c, x80, x81_c, x82, x84_c, x85_c, x86, x88, x92_c, x94_c, x96_c, x97_c, x99_c);
and (w737, x1_c, x2, x3, x4, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x11_c, x12, x13_c, x14, x15_c, x16, x17_c, x18_c, x19_c, x20, x21_c, x22_c, x23, x24_c, x25_c, x27_c, x28, x29, x30, x31_c, x32_c, x33, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50_c, x51_c, x52_c, x54, x55_c, x56_c, x57_c, x58_c, x59, x60_c, x61, x62, x64, x66_c, x67, x68, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76, x77, x78_c, x79, x81_c, x82_c, x83_c, x84, x85, x86_c, x87, x88, x89, x90_c, x91, x92_c, x93_c, x94_c, x95, x96, x97, x98_c, x99_c);
and (w738, x1, x3, x4, x6_c, x8_c, x11_c, x14, x15, x20_c, x22_c, x23, x24, x25, x26, x27_c, x30_c, x31_c, x33, x34_c, x35, x36_c, x37, x38, x39, x41_c, x43, x44_c, x48, x49_c, x50, x51, x53_c, x55_c, x56_c, x58, x59, x60_c, x62, x63, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x73_c, x74, x76, x78_c, x80_c, x82_c, x83, x84, x85, x86, x87_c, x89_c, x90_c, x91_c, x93_c, x96, x97_c);
and (w739, x1, x6, x14, x19_c, x26_c, x33_c, x48, x53, x59_c, x70, x76, x78_c, x83, x95_c);
and (w740, x1, x4_c, x7, x8_c, x11_c, x14, x15_c, x17, x18_c, x21_c, x22, x24, x25_c, x28_c, x31, x32, x34, x35, x38_c, x39_c, x41_c, x42, x48_c, x49, x50, x52, x57, x61_c, x62_c, x63_c, x64_c, x66_c, x67_c, x68_c, x69_c, x71_c, x73_c, x76, x77, x78_c, x80_c, x81, x82_c, x83, x84_c, x87_c, x93_c, x94, x97_c, x99);
and (w741, x2, x4, x10, x14_c, x19, x22, x24_c, x47, x55_c, x77, x79, x81, x83);
and (w742, x0, x1_c, x3, x5_c, x7, x10, x26_c, x27_c, x31, x33_c, x34_c, x39_c, x44_c, x50_c, x52, x53, x54_c, x57, x58, x65_c, x90_c, x92_c, x95_c, x96, x97);
and (w743, x1, x5_c, x16, x17, x19_c, x26_c, x30_c, x35_c, x37, x39, x40_c, x46, x48_c, x49_c, x52, x63_c, x72, x73, x74_c, x76_c, x79, x81_c, x83_c, x84_c, x89_c);
and (w744, x0, x4_c, x15_c, x22_c, x25_c, x31_c, x33_c, x34, x35_c, x48_c, x60, x61_c, x62, x64_c, x67, x69, x72, x73_c, x81_c, x83, x89, x90_c, x94_c, x95, x96_c);
and (w745, x0_c, x1_c, x4_c, x10_c, x11_c, x16, x20_c, x25_c, x34, x35, x36, x50, x54, x55, x59_c, x64_c, x69_c, x70_c, x71, x81, x86_c, x90_c, x91, x92, x93_c, x96_c);
and (w746, x0_c, x1, x2, x3_c, x5, x6_c, x7_c, x8, x10_c, x11_c, x12, x13, x14, x15_c, x16_c, x17, x18, x19, x20, x21_c, x22, x23, x25_c, x28_c, x29, x30_c, x31_c, x32_c, x33, x34, x36_c, x37, x38, x39_c, x40, x41, x42, x43_c, x44_c, x45_c, x46, x48, x49_c, x51, x53, x54_c, x55_c, x56, x58, x59, x60_c, x61_c, x62_c, x63_c, x64, x65, x66, x67_c, x68, x69, x70, x71_c, x72_c, x74_c, x77, x78_c, x79_c, x80, x81, x82_c, x83, x84_c, x85, x86, x87, x88_c, x89_c, x90, x91_c, x93, x95_c, x96, x97, x98_c);
and (w747, x0_c, x1_c, x3, x4, x5, x7, x8_c, x10_c, x13, x16_c, x18, x19, x20, x22, x24, x25_c, x26_c, x28_c, x29_c, x30, x33_c, x35, x36, x38, x39, x40, x41_c, x43, x44_c, x45_c, x46_c, x50_c, x52, x53_c, x54_c, x57, x58_c, x60_c, x61_c, x62, x64_c, x65, x68_c, x70, x71_c, x72, x73_c, x74, x75_c, x76, x81_c, x83_c, x85, x86, x87_c, x89, x94, x95_c, x96_c);
and (w748, x0_c, x4_c, x5_c, x6_c, x8_c, x9_c, x12_c, x13, x14_c, x16_c, x17, x18_c, x20_c, x22, x25_c, x26, x27, x29, x30_c, x31_c, x32_c, x36_c, x38, x39_c, x41_c, x43, x44, x45, x48_c, x49, x50_c, x51, x52, x53, x54, x55_c, x56_c, x57_c, x58_c, x60_c, x61, x62, x64, x65, x66, x68, x70, x71, x72_c, x74, x75_c, x76, x77, x78, x79_c, x81_c, x84_c, x85, x88_c, x89, x90, x91_c, x92_c, x97_c, x98_c, x99);
and (w749, x2_c, x3, x14, x15, x16, x19_c, x21_c, x22_c, x23, x24_c, x25_c, x27, x29_c, x30, x32_c, x33_c, x34, x35_c, x37, x39, x40_c, x42_c, x44_c, x47, x49_c, x55_c, x56, x60_c, x64, x66, x68_c, x69, x70, x72_c, x74_c, x76, x77_c, x78, x79_c, x82_c, x87, x88_c, x91, x92_c, x93, x95, x96, x97, x98, x99);
and (w750, x0_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8_c, x9_c, x10, x11, x12_c, x13, x14_c, x15_c, x16, x17, x19, x20_c, x21_c, x22_c, x23, x24_c, x25_c, x26, x27, x28, x29_c, x30, x31_c, x32_c, x33_c, x34_c, x35, x36, x37_c, x38, x39_c, x40, x41, x42, x43_c, x44_c, x45_c, x46_c, x47_c, x48_c, x49_c, x50_c, x51, x52, x53_c, x54_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63, x64_c, x65, x66_c, x67_c, x68_c, x69_c, x70_c, x71, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79, x80, x81, x82, x83_c, x85, x86, x87_c, x88, x89_c, x90, x92_c, x94, x95_c, x96_c, x97, x98, x99_c);
and (w751, x2, x5, x6_c, x7_c, x8, x12, x16, x17, x19_c, x21_c, x25_c, x27_c, x29_c, x30_c, x35, x36, x38_c, x39_c, x42_c, x47_c, x50, x51_c, x52_c, x53, x58_c, x59, x65_c, x70_c, x72_c, x73, x76_c, x78, x79, x81_c, x82_c, x83, x85_c, x90_c, x91_c, x93_c, x94, x95, x97, x99);
and (w752, x7, x17_c, x18, x19_c, x20_c, x23_c, x24_c, x29_c, x30, x33, x44, x48, x52, x55_c, x57_c, x58, x66, x67, x73_c, x76_c, x77_c, x79, x80_c, x85_c, x86_c, x87, x89, x95_c, x96_c, x97_c, x99);
and (w753, x0, x1, x2, x3, x5, x6_c, x7, x8, x9_c, x10_c, x11_c, x12_c, x13_c, x14, x15, x16, x18, x19, x20, x21, x22_c, x23, x24, x26, x27_c, x28_c, x29, x32_c, x33_c, x35_c, x36, x37, x38, x39_c, x41, x43, x44, x45_c, x46, x47_c, x48, x49_c, x52, x54, x56_c, x58, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66, x67_c, x68_c, x69_c, x70_c, x71, x72_c, x73, x74_c, x75_c, x76_c, x78_c, x79, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x88, x89_c, x90_c, x91, x92, x93_c, x94, x95, x96_c, x97, x99_c);
and (w754, x4_c, x6_c, x8, x10_c, x11, x13, x16_c, x18, x19_c, x22, x23_c, x24_c, x35, x38_c, x39_c, x41_c, x43, x46, x48, x49_c, x50, x54_c, x58_c, x63_c, x64_c, x68_c, x70, x73, x74_c, x76, x78_c, x80_c, x81_c, x84_c, x85, x87, x93_c, x95_c, x97_c, x98_c);
and (w755, x2_c, x3, x7, x11, x14, x16_c, x18_c, x19_c, x25, x38, x47_c, x48_c, x54_c, x55, x59, x60_c, x61_c, x67, x68, x69_c, x71_c, x72_c, x73, x75, x76_c, x79_c, x80, x84, x85_c, x87, x89_c, x90_c, x91, x93, x94, x95, x96_c, x98_c);
and (w756, x3_c, x4_c, x5, x7_c, x8_c, x9_c, x11, x14, x15_c, x17_c, x18_c, x21_c, x24, x32_c, x33, x35_c, x40_c, x41, x43_c, x44, x49, x52_c, x53, x59_c, x62, x63_c, x65, x66_c, x70_c, x72_c, x73, x78, x79_c, x82_c, x86, x89_c, x92_c, x93_c, x96, x97, x99);
and (w757, x0, x5_c, x10, x12, x18_c, x23, x24_c, x25_c, x27, x36, x37_c, x44, x49_c, x53_c, x64_c, x65, x78, x82, x87_c, x93, x95, x97_c, x98);
and (w758, x5_c, x10_c, x20_c, x32, x35, x36, x38, x40_c, x45, x46_c, x47_c, x51, x52_c, x63_c, x66, x73, x77, x79, x90, x91, x93);
and (w759, x1_c, x7_c, x8_c, x9_c, x13_c, x15_c, x17, x19, x20, x24, x25, x28, x31, x43_c, x44_c, x48, x49, x53, x54_c, x55_c, x60_c, x61, x62, x63_c, x64_c, x68_c, x72, x76_c, x79_c, x82, x85_c, x88, x89_c, x96_c);
and (w760, x0_c, x1_c, x2_c, x3, x4_c, x5, x6, x7_c, x8_c, x9, x10_c, x11_c, x12, x13, x14, x15_c, x16, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x24, x25_c, x26_c, x28_c, x29, x31, x32_c, x33, x34_c, x35, x36, x37_c, x38_c, x39_c, x41, x42, x43_c, x44, x45, x46, x47_c, x48, x49, x50_c, x51, x52, x53, x54, x55, x56, x57, x58, x59_c, x60_c, x61_c, x62_c, x63, x64, x65, x66_c, x68, x69, x70, x71_c, x72_c, x73_c, x74, x75, x76, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84, x85, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92_c, x93, x94_c, x95, x96, x97_c, x98, x99);
and (w761, x0, x1_c, x2_c, x3_c, x4, x5_c, x6, x7_c, x8, x9_c, x10, x11, x12_c, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x20, x21, x22_c, x23_c, x24, x25, x26_c, x27, x28, x29, x30, x31, x32, x33_c, x34_c, x35, x36, x37_c, x38, x39, x40, x41_c, x42, x43_c, x44, x45, x46_c, x47_c, x48_c, x49, x50, x51, x52_c, x53, x54, x55_c, x56, x57_c, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75, x76_c, x77, x78, x79, x80_c, x81, x82_c, x83, x84, x85_c, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93_c, x94, x95, x96, x97, x98_c, x99);
and (w762, x0, x1, x2, x3_c, x5_c, x6_c, x7_c, x8, x9_c, x10, x11, x12_c, x13, x14, x15_c, x16_c, x17_c, x20, x22_c, x23, x24_c, x25_c, x26_c, x27_c, x28, x29, x30_c, x31_c, x33, x34_c, x36_c, x37, x38_c, x39_c, x40_c, x41_c, x42_c, x43, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52_c, x53, x54, x57_c, x58, x59, x60, x61_c, x62, x63_c, x64_c, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73, x76, x77_c, x78_c, x79_c, x80, x81_c, x82, x83_c, x84, x86, x87, x88, x89, x90_c, x91, x92_c, x93, x94_c, x96_c, x97, x98_c, x99_c);
and (w763, x1, x4_c, x5_c, x6, x7_c, x8_c, x11, x12_c, x13_c, x15, x16, x20, x22, x26_c, x28, x30_c, x32_c, x34_c, x35_c, x36, x37_c, x43_c, x44, x45, x47_c, x49_c, x51, x53, x54_c, x56_c, x57, x58, x59_c, x60, x61, x62_c, x66_c, x67, x68, x72_c, x73_c, x78, x83, x84_c, x85, x86_c, x87_c, x88_c, x89_c, x92_c, x93_c, x96, x97, x99);
and (w764, x0_c, x3, x15_c, x16_c, x18_c, x23, x27, x33_c, x34_c, x38, x42, x43_c, x46_c, x47_c, x48_c, x51, x60, x61_c, x63, x64, x68_c, x70_c, x74_c, x79_c, x82_c, x84_c, x85_c, x86, x87, x88_c, x89_c, x90_c, x91, x99);
and (w765, x0, x1_c, x2, x3_c, x4_c, x5_c, x6_c, x7, x8, x9, x10_c, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17, x18, x19_c, x20, x21_c, x22, x23, x24, x25, x26, x27, x28, x29_c, x30_c, x31_c, x32, x33, x34, x35, x36, x37, x38_c, x39_c, x40, x41, x42, x43_c, x44, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51, x52, x53, x54, x55_c, x56_c, x57, x58, x59_c, x60_c, x61, x62_c, x63_c, x64_c, x65, x66_c, x67_c, x68, x69_c, x70, x71_c, x72, x73_c, x74_c, x75_c, x76, x77, x78_c, x79, x80, x81, x82, x83, x84_c, x85, x86_c, x87, x88, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98, x99);
and (w766, x6_c, x21_c, x39_c, x55_c, x57_c, x62, x65_c, x67, x72, x75, x95, x96);
and (w767, x0_c, x1_c, x2_c, x3, x5, x6, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14, x15, x17_c, x18, x20, x21, x22_c, x23_c, x24_c, x25, x28, x29, x31, x32_c, x33_c, x34, x35, x36, x37, x38, x39, x40, x41, x42_c, x43_c, x44_c, x45, x46_c, x47, x48_c, x49, x50_c, x51, x53, x54, x56, x58_c, x60_c, x61_c, x62_c, x63_c, x65_c, x66_c, x68, x69_c, x70_c, x71_c, x73_c, x74_c, x75, x76_c, x77_c, x78_c, x79, x82, x83_c, x84, x86, x87, x88, x89_c, x91, x93, x94_c, x95, x96_c, x97_c, x98, x99);
and (w768, x0, x3_c, x20_c, x22, x25_c, x28_c, x36, x37_c, x38_c, x46_c, x47, x49_c, x51, x54, x60, x61, x62_c, x75, x84_c, x85_c, x97_c);
and (w769, x0_c, x1_c, x2, x3_c, x5_c, x6_c, x7, x11_c, x12_c, x13, x15, x17_c, x18_c, x19_c, x20_c, x21_c, x25_c, x28_c, x33_c, x35, x37, x38_c, x39_c, x42_c, x44, x50, x51_c, x52_c, x53, x54_c, x56_c, x57, x58_c, x59, x60_c, x63, x64_c, x65, x66, x67_c, x68, x74_c, x76_c, x77, x78, x79_c, x82, x83, x84_c, x85, x88, x89, x90, x95_c, x96, x98_c, x99);
and (w770, x0_c, x2, x6, x9_c, x15, x17, x21_c, x22, x24, x26_c, x27, x29, x30_c, x32, x38_c, x40_c, x41, x44_c, x45, x47, x48, x49_c, x50, x52_c, x53, x54_c, x58_c, x60, x61_c, x64, x67, x69, x71_c, x72, x73, x74_c, x77, x78, x79_c, x87, x88_c, x89, x90, x91_c, x93, x95, x96_c);
and (w771, x0, x1_c, x2_c, x5_c, x6_c, x8, x16, x18, x24, x26_c, x28_c, x32, x35_c, x36, x38, x44, x45_c, x49_c, x50_c, x51, x56_c, x59_c, x62_c, x64_c, x65_c, x72, x73_c, x77, x80_c, x81_c, x82, x85_c, x87, x91_c, x92, x95_c, x96_c);
and (w772, x2_c, x11, x29_c);
and (w773, x0, x1, x2_c, x3_c, x4, x5, x6, x7_c, x8_c, x9, x10, x11_c, x12, x13, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21_c, x22, x23, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30, x31, x32, x33_c, x34, x35_c, x36_c, x37, x38, x39_c, x40_c, x41, x42, x43, x44_c, x45_c, x46, x47_c, x48, x49_c, x50_c, x51_c, x52_c, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61, x62_c, x63, x64, x65_c, x66, x67_c, x68_c, x69, x70, x71_c, x72_c, x73, x74, x75_c, x76, x77, x78, x79, x80, x81, x82_c, x83_c, x84, x85_c, x86_c, x87, x88_c, x89_c, x90, x91_c, x92, x93, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w774, x2, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10_c, x11_c, x12, x13, x14, x15_c, x16_c, x17_c, x18, x20_c, x21_c, x22_c, x23_c, x24, x25, x26, x27, x28, x29_c, x30_c, x31_c, x32_c, x33, x34_c, x35_c, x36, x38, x40, x42_c, x43, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x52_c, x53, x54, x55, x56, x57, x58_c, x59, x61_c, x62, x63, x64_c, x65, x66, x67, x69_c, x70, x71, x72, x75_c, x76_c, x77, x78_c, x79_c, x80, x81_c, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90_c, x91_c, x92, x93_c, x94, x95, x98_c, x99_c);
and (w775, x4_c, x7, x14, x16, x20_c, x25, x31, x32, x42_c, x50, x57_c, x65_c, x71, x74, x75_c, x80_c, x90);
and (w776, x1, x2_c, x6, x13_c, x14, x16_c, x17_c, x20, x21, x22, x24_c, x29_c, x31_c, x32, x34_c, x35_c, x38, x40_c, x41_c, x42_c, x47_c, x48, x49, x50_c, x52, x54, x56_c, x58_c, x60_c, x62_c, x64, x66, x70_c, x74, x76_c, x78, x79, x80_c, x83, x84, x85, x86_c, x91, x95_c);
and (w777, x0, x1, x2, x3_c, x4, x5_c, x6, x7_c, x8_c, x9_c, x10, x11_c, x12, x13, x14, x15_c, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24_c, x25, x26_c, x27, x28_c, x29_c, x30, x31_c, x32, x33_c, x34, x35, x36_c, x37_c, x38, x39, x40_c, x41, x42_c, x43, x44_c, x45_c, x46_c, x47_c, x48_c, x49, x50_c, x51, x52_c, x53_c, x54, x55, x56, x57, x58_c, x59, x60, x61, x62, x63, x64, x65, x66, x67_c, x68_c, x69_c, x70_c, x71, x72, x73, x74_c, x76, x77_c, x78_c, x79_c, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91, x92_c, x93_c, x94, x95, x96, x97_c, x98, x99);
and (w778, x19, x26_c, x34, x35, x38_c, x40, x44, x59, x60, x68, x78, x86_c, x87_c, x99_c);
and (w779, x0, x1, x2, x3, x5_c, x6_c, x7_c, x8_c, x9, x12_c, x13, x14, x15_c, x16, x17, x18, x20, x21, x24, x25_c, x28_c, x29, x30_c, x31, x32_c, x33, x34_c, x37, x38_c, x39_c, x40, x41, x43_c, x44_c, x45_c, x47, x48, x49_c, x52, x54_c, x57_c, x58_c, x59, x60, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68, x69, x70, x71_c, x73_c, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82, x83_c, x84_c, x85_c, x88, x90, x91, x92_c, x93_c, x94, x99_c);
and (w780, x0, x1, x2, x3, x4_c, x5, x8_c, x9_c, x10_c, x11_c, x12, x13, x14_c, x15, x16_c, x17_c, x18, x19_c, x20_c, x21, x22_c, x23, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32, x33, x34, x35, x36_c, x38_c, x39, x40_c, x41, x42, x44, x45_c, x46, x47, x48, x49, x52_c, x53_c, x55, x57_c, x59_c, x61_c, x62, x63, x64_c, x65_c, x66_c, x69_c, x70, x71, x72_c, x74, x75, x76_c, x77, x79, x81, x82, x83_c, x84, x86_c, x87, x88_c, x89_c, x91_c, x92, x94_c, x95_c, x96, x97_c, x98, x99_c);
and (w781, x0, x4, x5, x7, x9_c, x10, x14, x16, x17, x23, x24_c, x25_c, x32_c, x33_c, x40, x41, x46_c, x48, x51, x55_c, x58, x63_c, x70, x75, x79, x80_c, x85_c, x87_c, x88, x91, x94, x96);
and (w782, x1, x4, x7, x8_c, x11, x12, x13, x14, x19_c, x21, x22_c, x24, x27, x28_c, x38, x43_c, x53_c, x54, x55_c, x56_c, x59_c, x69_c, x72_c, x73_c, x74, x77, x83_c, x84, x85_c, x96_c, x98_c);
and (w783, x22_c, x24_c, x33_c, x37, x43_c, x53, x63, x65, x76, x90_c, x92_c, x96, x99);
and (w784, x0_c, x1_c, x2_c, x3, x4_c, x5, x6, x7, x8_c, x9, x10, x11, x12_c, x13_c, x14_c, x15, x16, x17, x18, x19_c, x20, x21_c, x22_c, x23, x24, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31, x32_c, x33, x34, x35_c, x36, x37, x38_c, x39_c, x40_c, x41, x42, x43_c, x44, x46, x47, x48, x49, x50_c, x51, x53_c, x54, x55_c, x56_c, x57, x58_c, x59, x60_c, x61_c, x62, x63_c, x64_c, x66, x67, x68, x69_c, x70, x71, x72, x73_c, x74_c, x75, x76, x77, x78, x79_c, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x86_c, x87_c, x88_c, x89_c, x90, x91, x92, x93, x94_c, x95, x96, x97_c, x98_c);
and (w785, x0, x1_c, x3, x4, x5, x6_c, x8_c, x9_c, x10, x12, x13_c, x14_c, x15_c, x16, x17_c, x18_c, x20, x21_c, x22, x24_c, x25, x26, x27, x28_c, x29, x30, x32, x33_c, x34_c, x36_c, x37, x39_c, x40, x41, x42, x43, x44, x45, x46, x47, x49_c, x50_c, x52_c, x55, x57_c, x58, x59_c, x60, x62_c, x63, x64, x65, x68_c, x70, x71, x72_c, x73, x75, x76_c, x78, x79_c, x80, x82_c, x83, x86, x87_c, x88, x89_c, x90, x91, x93_c, x94, x95, x97, x99_c);
and (w786, x0, x2, x7_c, x8_c, x11, x13_c, x18_c, x21_c, x27_c, x30_c, x31, x32, x40_c, x46, x47_c, x56_c, x67_c, x79_c, x80_c, x87, x88, x91, x93_c, x97, x98_c);
and (w787, x0_c, x1, x2, x3, x7, x8, x9_c, x10_c, x11, x12, x13_c, x14_c, x15, x17, x18, x20, x21_c, x22, x23_c, x24_c, x25, x26_c, x27, x29_c, x30_c, x31_c, x32, x33_c, x35, x36, x37_c, x39, x40_c, x41_c, x42_c, x43, x44, x47_c, x48_c, x49, x50, x52, x53, x54, x56_c, x57, x58_c, x59, x60, x61, x63_c, x64_c, x65, x66_c, x68_c, x69, x70, x72_c, x73, x74_c, x76, x77_c, x79, x80, x81, x85, x86, x87, x88, x89, x91_c, x92, x95_c, x96, x97, x99);
and (w788, x0, x1, x2_c, x3, x4_c, x5, x6, x7_c, x8_c, x10_c, x12_c, x14_c, x17, x18_c, x20_c, x21_c, x22_c, x24, x27, x28, x29_c, x31_c, x32_c, x35, x36, x37, x38_c, x39, x41_c, x42, x43_c, x44_c, x45, x47, x49_c, x50_c, x51_c, x53, x54, x56, x57, x58_c, x59, x60_c, x62_c, x65_c, x66, x68, x69_c, x70, x71_c, x72, x73, x74_c, x76, x77_c, x81_c, x83, x84, x85_c, x86, x87_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98_c);
and (w789, x0, x4, x31, x36, x41, x47_c, x54_c, x77_c, x80, x84_c, x87_c, x95_c, x96_c);
and (w790, x0_c, x1, x2_c, x3_c, x4, x5_c, x6, x7, x8, x9, x10_c, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x21, x22, x23_c, x24, x26, x27_c, x28, x29, x30_c, x31, x32, x33, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x43_c, x45_c, x46_c, x47_c, x48, x49_c, x50_c, x51, x52, x53, x54_c, x55_c, x56, x58_c, x59_c, x60_c, x61, x62_c, x63, x64, x65_c, x66, x67_c, x68, x69, x70, x71_c, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79_c, x81_c, x82, x83_c, x84_c, x85_c, x86, x87, x88, x89, x90_c, x91_c, x92, x93_c, x94, x95_c, x96, x97_c, x98_c, x99);
and (w791, x11, x12_c, x15, x17_c, x23_c, x27, x29_c, x31, x41_c, x46, x47_c, x54_c, x55, x60_c, x64, x70, x71, x73_c, x78, x86, x93_c, x95_c, x97);
and (w792, x0, x1, x3_c, x4, x7, x8_c, x9_c, x10_c, x11, x12_c, x14_c, x15_c, x16_c, x17_c, x18, x19, x21, x22_c, x25_c, x27_c, x29, x30_c, x31_c, x32, x33_c, x34, x35_c, x36, x37_c, x38_c, x39, x40_c, x41, x42_c, x43_c, x45_c, x46_c, x47_c, x48, x49, x50, x52, x53_c, x55, x56_c, x57, x58_c, x59, x60_c, x61, x62, x64, x65, x66, x67, x68_c, x70_c, x72, x73_c, x74_c, x75, x76_c, x77, x78_c, x79, x80_c, x81_c, x82_c, x83, x84_c, x85, x86_c, x87, x89, x90, x91, x93, x95_c, x96_c, x97_c, x98, x99);
and (w793, x0_c, x1_c, x2_c, x4, x6, x7, x8_c, x9, x11_c, x13_c, x17, x18, x19, x20, x22, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x35_c, x36, x38, x39, x41_c, x42_c, x43_c, x44, x45, x46_c, x47_c, x48_c, x49, x50_c, x53, x54, x55, x56_c, x57_c, x58, x60_c, x62, x65_c, x67, x68, x69, x72, x74_c, x76_c, x78, x79, x81, x82_c, x84, x85, x86_c, x87_c, x88_c, x90_c, x91, x92, x94, x95_c, x96_c, x99);
and (w794, x0, x1_c, x3, x5_c, x6, x7_c, x8_c, x10, x11, x12_c, x13, x14_c, x15_c, x16_c, x17_c, x19_c, x20, x22, x23_c, x24, x25_c, x26_c, x27, x29_c, x30_c, x31_c, x32, x33, x36_c, x39, x40, x41, x42, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x52_c, x53, x54, x55_c, x57_c, x58_c, x59, x60, x61_c, x63, x65_c, x66_c, x67_c, x68_c, x69_c, x70, x71, x72, x73_c, x74_c, x75, x77_c, x78_c, x79, x80_c, x82, x83, x84, x85_c, x87_c, x88, x89_c, x90_c, x91, x92_c, x93, x94_c, x96_c, x97, x98, x99);
and (w795, x4, x5_c, x9_c, x26_c, x35_c, x37, x42, x45, x49, x80, x84);
and (w796, x0, x1, x3, x6, x7_c, x9, x10, x11_c, x12_c, x13, x14_c, x15_c, x16_c, x17_c, x18, x19, x21_c, x23, x24_c, x25, x26, x27_c, x28, x30_c, x32, x33, x34_c, x36_c, x37, x40, x41_c, x43, x44, x45_c, x46, x47, x49_c, x51_c, x53, x54, x55, x56, x57, x59_c, x60_c, x62, x63_c, x65, x67_c, x68, x70_c, x71, x73, x75_c, x76, x77, x79, x81_c, x82, x83_c, x85, x86, x87, x88, x89_c, x91, x92, x94, x96, x98, x99_c);
and (w797, x0_c, x1, x2_c, x4, x5_c, x6_c, x8, x9_c, x10, x11, x12, x13, x16, x17, x18_c, x19, x21, x22_c, x23, x24_c, x25_c, x26, x30_c, x31, x32, x34_c, x35, x39, x42, x44, x46_c, x47_c, x48, x49_c, x51, x52_c, x53, x54, x56, x57_c, x58_c, x59_c, x61, x63, x64, x66, x67, x68, x72_c, x73, x74, x75, x77_c, x79, x80_c, x81, x82, x83, x84, x85_c, x86, x87_c, x88_c, x89_c, x90, x92, x94, x97, x98_c, x99_c);
and (w798, x53_c, x83_c);
and (w799, x0, x2, x7_c, x8, x11_c, x13, x14_c, x27, x28, x30, x53, x55_c, x63, x65, x81, x95, x98_c);
and (w800, x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x8_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16_c, x19, x20, x21_c, x22, x23, x24_c, x25_c, x27, x28, x29, x30, x32, x33_c, x34, x35_c, x36, x37, x38_c, x39, x40, x41_c, x42, x43, x44_c, x45, x46, x47_c, x48_c, x49_c, x50_c, x51, x52_c, x53, x54, x55_c, x56, x57_c, x58, x59_c, x60, x61_c, x62, x63_c, x64, x66_c, x67_c, x69, x70_c, x71_c, x73_c, x74, x76_c, x77_c, x78, x79, x80, x81_c, x82_c, x83, x84_c, x85_c, x86, x87, x88_c, x89_c, x90, x91, x92_c, x93_c, x94_c, x95_c, x96, x97_c, x98, x99_c);
and (w801, x0, x1, x2_c, x3, x4, x6_c, x7_c, x8, x9, x10, x11_c, x12_c, x13, x14, x15, x17_c, x18_c, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28, x29_c, x30_c, x31_c, x32, x33_c, x36_c, x37_c, x38, x39_c, x40_c, x42_c, x43_c, x44, x45, x46_c, x47, x48_c, x49, x50, x51_c, x52, x53, x54, x55, x57_c, x58_c, x59, x60_c, x61, x62, x63, x64_c, x65, x66_c, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80, x81, x82_c, x83_c, x84_c, x85, x86, x87_c, x88, x89, x90, x91, x92, x93_c, x94, x95, x96, x98_c, x99_c);
and (w802, x0, x1_c, x3, x4_c, x5_c, x6, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x15, x16, x17, x18, x20_c, x21_c, x22_c, x23_c, x25_c, x28, x29, x30, x31_c, x36_c, x37_c, x38_c, x39_c, x40, x41, x42, x44, x46_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55_c, x58, x61_c, x62_c, x64, x65_c, x66, x67, x69_c, x70, x72_c, x73_c, x74_c, x75_c, x76, x78_c, x79_c, x80, x81, x82, x84, x85_c, x86_c, x87_c, x88_c, x91, x92_c, x94, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w803, x0, x1, x2_c, x4, x5, x6, x8_c, x9, x11_c, x12_c, x13_c, x14, x17, x27_c, x29, x31, x34, x36_c, x38_c, x41, x44, x45, x48_c, x49, x50_c, x51, x52_c, x59, x63_c, x64_c, x69, x70_c, x71, x74_c, x75, x80, x83, x84_c, x85, x87, x89, x92, x97, x98, x99);
and (w804, x20_c, x21, x35, x40, x54_c, x70_c, x74_c, x90);
and (w805, x0, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9_c, x10, x11_c, x12, x13_c, x14, x15, x16_c, x17_c, x18, x19_c, x20_c, x22, x23_c, x24_c, x25_c, x26_c, x27_c, x28, x29, x30_c, x31, x33_c, x34_c, x35_c, x36_c, x37_c, x38_c, x39_c, x40, x41_c, x42, x43_c, x44_c, x45, x46_c, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x55, x56_c, x57_c, x58, x59_c, x60, x61, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x72_c, x73, x74, x75_c, x76, x77, x78_c, x79, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88_c, x89, x90, x91, x92_c, x93, x96_c, x97, x98, x99);
and (w806, x0_c, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x8_c, x9, x10, x11, x12, x13_c, x14_c, x15_c, x16, x17, x18_c, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33, x34, x35_c, x36_c, x37_c, x38, x39, x40_c, x41_c, x42_c, x43_c, x45, x46, x47_c, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66, x67_c, x68, x69_c, x70_c, x71, x72_c, x73, x74, x75, x76, x77_c, x78_c, x79, x80, x81_c, x82_c, x83_c, x84, x85_c, x86, x87, x88_c, x89_c, x90, x91_c, x92, x93, x94_c, x95_c, x96_c, x97_c, x98_c, x99_c);
and (w807, x0, x1_c, x2_c, x3_c, x4_c, x5, x6_c, x7, x8_c, x9, x10_c, x11_c, x12, x13, x14_c, x15_c, x16, x17_c, x18_c, x19, x20, x21_c, x22_c, x23_c, x24, x25, x26, x27_c, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34_c, x35, x36_c, x37, x38, x39, x40, x41_c, x42_c, x43, x44_c, x45_c, x46_c, x47, x49, x50_c, x51, x52_c, x54, x56_c, x57_c, x58_c, x59, x60_c, x61, x62, x63_c, x65, x66_c, x67_c, x68, x69_c, x70, x71, x72, x73_c, x74, x75_c, x76_c, x77, x78, x79_c, x81, x82_c, x83, x84_c, x85_c, x86, x87_c, x88_c, x90, x91, x92_c, x93_c, x94, x95, x96, x97, x98, x99_c);
and (w808, x1, x5, x12_c, x19_c, x30, x38_c, x45_c, x47, x48, x49_c, x50, x52_c, x54, x57_c, x60, x73_c, x77, x80_c, x82_c, x88, x96, x97);
and (w809, x3_c, x9_c, x15_c, x18_c, x19_c, x24_c, x26, x28, x29_c, x30, x31, x33_c, x36, x39_c, x41, x42_c, x43, x45, x49, x56_c, x57_c, x58_c, x59_c, x61, x62, x63_c, x71_c, x74, x77_c, x80, x81_c, x82, x83_c, x91_c, x93_c, x94_c, x95, x97, x98_c);
and (w810, x0, x1, x2_c, x3, x4, x5_c, x6_c, x7, x8, x9_c, x10_c, x11, x12_c, x13, x14, x15, x16_c, x17, x18_c, x19, x21_c, x22, x23_c, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34_c, x35, x36, x38, x39_c, x40_c, x41, x42_c, x43_c, x44_c, x45_c, x46_c, x47, x48, x49_c, x50, x51, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60_c, x61_c, x62, x63, x64, x65, x66, x67_c, x68_c, x69, x70, x71, x72, x73, x74, x75_c, x76, x77, x78_c, x79_c, x80_c, x81, x82_c, x83, x84_c, x85, x86_c, x87_c, x88, x89, x90_c, x91_c, x92, x93, x94, x95, x96, x97, x98_c, x99_c);
and (w811, x15_c, x19, x23_c, x35_c, x60, x84, x88_c);
and (w812, x2, x6, x8, x11_c, x12_c, x13, x18, x26, x36_c, x42, x43_c, x50, x52_c, x57_c, x61_c, x67, x70, x72_c, x78, x80_c, x82, x86, x88_c, x89_c, x90_c, x95, x97, x99_c);
and (w813, x0_c, x1_c, x2, x3_c, x4_c, x5, x6_c, x8_c, x9_c, x10_c, x11, x12_c, x13_c, x14, x15_c, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29, x30_c, x31_c, x32, x33_c, x34_c, x36_c, x37_c, x38, x39, x40_c, x41, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48, x49_c, x50_c, x51_c, x52, x53_c, x54, x55_c, x56_c, x57_c, x58, x59_c, x60, x61_c, x62, x63_c, x64_c, x65_c, x66_c, x67, x68, x69_c, x70_c, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78_c, x79_c, x80, x81, x82, x83_c, x84_c, x85, x86, x87_c, x88_c, x89_c, x90_c, x91_c, x92_c, x93_c, x94, x95_c, x96_c, x97, x98_c, x99);
and (w814, x2, x3_c, x4_c, x5_c, x7_c, x8_c, x9, x10, x11, x12, x13_c, x14, x15_c, x16, x17_c, x18, x19_c, x20_c, x24_c, x25, x26_c, x27_c, x28_c, x29, x30, x31, x33_c, x34_c, x35, x36_c, x37_c, x38_c, x39_c, x40_c, x41_c, x42, x43_c, x44_c, x45, x46, x47, x49, x50_c, x52, x54_c, x55_c, x56, x57_c, x58, x59_c, x60_c, x61_c, x62_c, x63_c, x64_c, x65, x66, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x78_c, x79, x80_c, x82, x85_c, x86, x87, x88_c, x89_c, x90_c, x93_c, x94_c, x95, x96, x97, x98_c, x99_c);
and (w815, x0_c, x1, x2, x3, x4, x6_c, x7, x8_c, x9_c, x10_c, x11_c, x12, x13_c, x14_c, x15_c, x17, x18, x20_c, x21_c, x22_c, x23, x24, x25_c, x26, x27, x28_c, x29, x30_c, x31, x32, x33, x34, x36, x37, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46_c, x48, x49, x50, x51_c, x52_c, x53, x55_c, x56_c, x57, x58, x59, x61_c, x63, x64_c, x65_c, x66_c, x67_c, x68, x69_c, x70_c, x71_c, x73, x75, x78_c, x80, x81_c, x82, x83_c, x84_c, x85_c, x86_c, x87, x88, x89, x90, x91, x92, x93_c, x94, x96_c, x98, x99);
and (w816, x0, x2_c, x6_c, x8_c, x9_c, x10_c, x11_c, x13, x16_c, x19, x20_c, x23_c, x24_c, x25_c, x26_c, x29_c, x30, x31, x33, x36, x39_c, x40_c, x41, x48_c, x50_c, x53_c, x56_c, x57_c, x58, x59, x60, x61_c, x64_c, x65, x71, x77, x78_c, x81, x83, x86, x87, x89_c, x90, x91, x93, x96_c, x98, x99);
and (w817, x0, x1, x2, x3, x4, x6, x7, x8, x9, x10, x11_c, x12_c, x13, x14_c, x15_c, x16, x18, x19_c, x20_c, x22, x23_c, x24, x25, x26_c, x27, x28, x29, x30, x31_c, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38_c, x39_c, x40_c, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49, x50_c, x51_c, x52, x53, x54, x56, x57_c, x58, x60_c, x61_c, x62, x63_c, x64_c, x65_c, x66, x67_c, x68, x69, x70_c, x72, x73_c, x74, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x82, x83_c, x84_c, x85_c, x86_c, x87, x88, x89, x90, x91_c, x92_c, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w818, x0_c, x1, x2_c, x3_c, x4, x5_c, x6, x7_c, x9_c, x10, x11, x12_c, x13_c, x14, x15_c, x16_c, x17, x18_c, x19_c, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x29, x30, x31, x32, x33, x34_c, x35_c, x36_c, x37, x38_c, x39_c, x40, x41, x42_c, x43, x44, x46_c, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54_c, x55, x57_c, x58_c, x59_c, x60, x61_c, x62_c, x63, x64_c, x65, x67_c, x68_c, x69_c, x70, x71, x72, x73_c, x74, x75_c, x76, x77, x78, x79, x80, x81_c, x82, x83_c, x84_c, x85_c, x86_c, x87_c, x88, x89_c, x90, x91_c, x92_c, x93, x94_c, x95_c, x97, x99_c);
and (w819, x2_c, x3, x5, x6, x7, x8, x9_c, x10_c, x12, x13, x14_c, x16_c, x21, x24_c, x27_c, x29_c, x30, x32, x34, x35, x38, x40, x42, x44_c, x45, x48, x49, x50_c, x51_c, x52, x53, x55, x56, x59, x61, x62, x63, x67_c, x68, x70, x74, x78, x83, x84_c, x86_c, x88_c, x89_c, x91, x96, x97, x98_c);
and (w820, x0, x2, x4_c, x5_c, x7_c, x8_c, x10_c, x11, x12, x13, x14, x16, x18, x19_c, x20_c, x22_c, x24, x31_c, x32_c, x33, x34_c, x38, x39_c, x40_c, x42_c, x43, x47_c, x48_c, x49, x51, x52_c, x53_c, x54, x57, x59_c, x60, x63, x64_c, x66_c, x67_c, x68_c, x69, x70_c, x71, x72, x74_c, x76_c, x77, x78, x80, x82, x84_c, x86_c, x87, x88_c, x95, x96_c);
and (w821, x0, x1_c, x2_c, x4, x10_c, x16_c, x17, x18_c, x19, x22, x24_c, x27, x31_c, x32, x35, x36_c, x39, x45, x46, x47_c, x50, x53_c, x54, x59_c, x60, x61, x64, x66_c, x72, x74, x78_c, x86, x91_c, x92_c, x95, x97_c);
and (w822, x23, x62, x66_c, x67, x70_c);
and (w823, x1, x3_c, x11_c, x13_c, x19, x20, x25, x26_c, x27, x32_c, x34_c, x41_c, x43_c, x44_c, x45, x53, x57, x59, x61, x70, x83, x88, x94, x96, x97_c);
and (w824, x0, x2, x8, x9_c, x10, x13_c, x15_c, x18, x19, x20_c, x21, x23, x24, x25_c, x27, x32, x34, x35, x36_c, x39, x45_c, x49_c, x50, x52, x53_c, x55, x62_c, x64_c, x65, x67_c, x68, x70, x73, x74_c, x75_c, x79_c, x81, x82_c, x83_c, x85_c, x86_c, x88, x92_c, x94_c, x96, x98);
and (w825, x3_c, x4, x5, x6_c, x8_c, x10_c, x12, x14, x15_c, x17_c, x19_c, x20, x21, x24, x29_c, x32_c, x33_c, x34, x36, x40_c, x48_c, x50_c, x55_c, x56, x60, x61_c, x62, x66, x68, x72_c, x73, x76, x78_c, x79_c, x84_c, x87, x90, x92_c);
and (w826, x0, x1_c, x2_c, x3, x5_c, x6_c, x7_c, x8_c, x11, x12_c, x13, x17_c, x19_c, x20, x23_c, x24_c, x25_c, x26, x28, x30, x31, x33_c, x34_c, x35, x36, x37, x38_c, x39_c, x41, x42, x43, x44, x45_c, x46, x47_c, x48, x49_c, x52_c, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61_c, x62, x64, x65_c, x68_c, x70_c, x71_c, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80_c, x82_c, x83, x84, x85, x87_c, x88_c, x89, x90, x91_c, x93_c, x94, x95, x96_c, x97_c, x99_c);
and (w827, x13, x20_c, x21, x26, x30_c, x31, x36, x39, x40, x43, x44_c, x47, x59_c, x68, x71_c, x76, x80, x81, x86_c, x87, x88_c, x99);
and (w828, x15_c, x19, x23_c, x35, x45, x46, x60_c, x63, x69_c, x72, x79, x84, x90_c, x93);
and (w829, x14, x17, x22, x25_c, x33, x39_c, x45, x63, x69, x77_c, x83_c, x84_c, x97_c);
and (w830, x1, x3, x5, x6_c, x7_c, x9_c, x12, x16_c, x20, x21_c, x22, x24_c, x28_c, x29, x34_c, x42_c, x45, x46_c, x54_c, x57_c, x58_c, x63, x69, x70, x73, x78_c, x83, x84_c, x88_c, x89, x96_c, x98_c, x99_c);
and (w831, x0, x1, x3, x4_c, x5, x6, x7, x8_c, x9_c, x10_c, x12_c, x13_c, x14_c, x15, x16_c, x17_c, x19, x21, x22_c, x23_c, x24, x27, x28_c, x29, x30_c, x31_c, x32, x33, x34, x35_c, x36, x38, x39_c, x41_c, x42, x43, x44_c, x45_c, x46, x47, x48_c, x51, x52, x53_c, x54_c, x55, x56, x58, x60_c, x61_c, x63, x64_c, x65, x66, x67_c, x68, x69, x70, x72_c, x73, x74_c, x75_c, x76, x77, x79, x80, x82, x83, x84_c, x85, x89_c, x90_c, x91_c, x93_c, x94_c, x95_c, x97_c, x99);
and (w832, x1_c, x2, x5, x6, x8_c, x9, x10_c, x15, x16_c, x23_c, x27, x28, x29, x31_c, x40, x41_c, x43_c, x44, x46, x48_c, x52, x53, x54, x56_c, x57, x60_c, x61, x62, x63, x67, x68, x82_c, x88_c, x90_c, x92, x93_c, x98_c);
and (w833, x0, x1, x2_c, x3_c, x4, x5_c, x6_c, x7_c, x8_c, x9, x11_c, x12, x13, x14_c, x15, x16, x17, x18_c, x19, x20_c, x21_c, x22_c, x23_c, x24, x25_c, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33_c, x34_c, x35, x36, x37, x38, x39_c, x40, x41, x42, x43, x44_c, x45_c, x46, x47_c, x48, x49_c, x50_c, x51, x52_c, x53, x54_c, x55_c, x56, x57, x58, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66_c, x67_c, x68_c, x69, x70, x71, x72_c, x73, x74, x75_c, x76_c, x77, x78, x79, x80, x81, x82_c, x83_c, x84, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91, x92, x93, x94, x95, x96_c, x97_c, x98_c, x99);
and (w834, x0_c, x1, x3, x4_c, x5, x6, x7_c, x8_c, x10, x11_c, x12_c, x14, x15_c, x16_c, x17, x18, x20_c, x21_c, x22_c, x23_c, x24, x25, x26_c, x27_c, x28_c, x29, x30, x31_c, x32, x33_c, x34_c, x36_c, x38, x39_c, x40_c, x41, x43, x44_c, x46, x47_c, x48_c, x50, x51_c, x52, x53_c, x54_c, x55_c, x56_c, x57, x58, x60, x61_c, x62, x63_c, x64_c, x65, x66, x67_c, x70_c, x71, x72, x73_c, x75, x76_c, x79_c, x80_c, x81_c, x82, x83_c, x84_c, x85, x86, x87_c, x88, x92_c, x93, x94_c, x95_c, x96, x97_c, x98, x99);
and (w835, x2_c, x4_c, x8, x9, x11, x12, x16_c, x19_c, x21_c, x23_c, x25, x27_c, x28_c, x30_c, x31, x33, x34_c, x36_c, x37, x38_c, x41, x42, x45, x47, x50_c, x51_c, x52, x53_c, x56_c, x58, x62, x63_c, x64, x65_c, x67_c, x69_c, x72, x74, x76, x79_c, x80_c, x81_c, x83, x85, x87, x92, x96_c, x98_c);
and (w836, x0, x3, x5_c, x6_c, x7_c, x9, x13, x15, x16, x20, x21_c, x24, x26_c, x27, x28, x30_c, x31, x32_c, x33_c, x35, x36, x37_c, x38, x41, x42, x43_c, x45, x46, x48_c, x49, x52, x53, x54, x56, x57_c, x58, x60_c, x61, x62_c, x64, x66, x67_c, x68_c, x70_c, x71, x72_c, x73, x75_c, x76_c, x78_c, x83, x86, x87_c, x89_c, x94, x99_c);
and (w837, x7, x12, x14_c, x18, x20, x28_c, x35_c, x36_c, x38, x43, x55_c, x63_c, x74_c, x80, x85_c, x87, x89_c, x91, x92, x94, x95);
and (w838, x3, x5_c, x8, x14_c, x15, x30_c, x35, x36, x38, x39, x40, x49, x61, x62_c, x76_c);
and (w839, x8_c, x37, x54);
and (w840, x1, x2, x4, x15_c, x18_c, x19_c, x21, x26_c, x28_c, x29_c, x38, x39_c, x47_c, x48, x49_c, x53_c, x58, x59, x62_c, x77, x79, x80, x82_c, x86_c, x87);
and (w841, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8, x9, x13, x14, x15_c, x17_c, x18_c, x19, x21, x22_c, x23_c, x24, x25_c, x26, x27_c, x28_c, x29_c, x31_c, x33_c, x35, x36_c, x38, x39_c, x40_c, x42_c, x43, x46_c, x47, x48, x49, x50_c, x51, x52, x53_c, x54_c, x55, x56, x57, x58, x59_c, x60_c, x61_c, x63_c, x64, x66, x67, x68, x69_c, x70, x71_c, x72_c, x73_c, x74, x75, x77_c, x78_c, x83, x85_c, x86, x88, x90, x91_c, x93_c, x95, x96, x97_c, x98, x99_c);
and (w842, x1_c, x4_c, x8_c, x9_c, x10, x13_c, x14_c, x18, x23, x30_c, x33, x38, x39, x40, x42, x44_c, x50, x51_c, x56_c, x57, x58_c, x76, x84_c, x91, x94, x95_c, x98, x99);
and (w843, x1_c, x2, x4_c, x5, x7_c, x9, x11_c, x14_c, x15, x17, x18_c, x20_c, x21_c, x22_c, x23_c, x25, x26_c, x28, x29, x30, x31_c, x32, x33_c, x34, x36, x38, x39_c, x40, x43_c, x44_c, x47_c, x48_c, x50, x54, x58_c, x60_c, x61_c, x62, x64, x66_c, x68, x71, x73, x74, x75, x79, x81_c, x82_c, x84, x85, x88_c, x90_c, x91, x92_c, x98);
and (w844, x1_c, x2_c, x3, x4, x5, x11_c, x13, x14_c, x17, x18_c, x23, x24_c, x25_c, x27, x28, x31_c, x32_c, x33_c, x34_c, x38, x40, x42, x43_c, x44_c, x45, x48_c, x51, x52, x53_c, x54, x56, x57_c, x59_c, x62, x66, x67, x69, x73, x81, x82_c, x87, x90_c, x91_c, x92, x94_c, x97, x98, x99);
and (w845, x2_c, x3_c, x6, x8_c, x11_c, x13_c, x16, x18, x19_c, x24, x25, x26_c, x29_c, x33_c, x34, x35_c, x36, x38_c, x39_c, x40, x44, x45_c, x51, x52_c, x59, x61_c, x67, x76, x80_c, x81, x82_c, x84_c, x85, x86_c, x88, x89_c, x96, x97_c, x98_c);
and (w846, x0_c, x2_c, x4, x5, x7, x8_c, x9, x10_c, x12, x13_c, x20_c, x21, x24, x25, x29, x31_c, x32, x33, x34, x35, x36, x37_c, x38, x45, x49, x50_c, x54, x55_c, x56, x58_c, x59, x62_c, x63_c, x65_c, x73_c, x75_c, x77, x79, x80_c, x81, x83, x86_c, x90_c, x91_c, x92_c, x93, x94_c, x97_c, x98, x99_c);
and (w847, x2_c, x5_c, x7, x8_c, x12, x15_c, x16, x18_c, x21, x22_c, x23_c, x24, x26_c, x30, x33, x38_c, x40, x45_c, x47_c, x54_c, x55, x56, x57_c, x60, x63_c, x64, x65, x67, x68_c, x69_c, x70_c, x75_c, x78_c, x79, x80_c, x83_c, x87, x88_c, x90, x92_c, x98);
and (w848, x1, x4, x5_c, x6_c, x8_c, x11, x12, x13, x14_c, x15_c, x16, x18, x19, x20, x21_c, x23, x24_c, x25_c, x27, x28_c, x29, x30_c, x35_c, x37_c, x40_c, x41, x42_c, x46_c, x48, x49, x51_c, x52_c, x53, x54, x55_c, x56_c, x57, x58, x59_c, x60_c, x61_c, x62_c, x66_c, x67_c, x68, x69_c, x70, x71_c, x72, x73_c, x74, x76, x77, x78_c, x79, x80_c, x82_c, x83, x84, x85, x86_c, x87_c, x91_c, x92_c, x93, x94, x96, x97_c, x98_c, x99);
and (w849, x1, x14_c, x26_c);
and (w850, x4_c, x5, x7_c, x12, x14, x15, x21_c, x23_c, x30_c, x31, x36_c, x37_c, x41_c, x45_c, x49, x51, x52, x54_c, x55, x61, x62_c, x66_c, x70, x75_c, x77_c, x90_c, x92, x96);
and (w851, x6_c, x17, x25_c, x38, x48_c, x58_c, x66_c, x68_c);
and (w852, x0, x1, x2_c, x3_c, x4, x5_c, x9_c, x10, x11_c, x12, x13_c, x14, x15, x17, x18, x19, x21, x23, x24, x25, x26, x27_c, x28_c, x32_c, x33_c, x34_c, x36_c, x38_c, x39, x40, x41_c, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x50_c, x51, x52, x55_c, x57_c, x58_c, x59_c, x63_c, x64, x65, x66_c, x69, x70_c, x75, x76_c, x77, x78_c, x83, x85, x86, x87, x88, x89, x91_c, x92, x93, x94_c, x95, x96, x97, x98, x99_c);
and (w853, x2_c, x3_c, x4, x6, x7, x8, x9_c, x10, x11, x12_c, x13, x16, x17_c, x18_c, x19_c, x21_c, x22, x24_c, x25, x26, x28_c, x29, x30, x31_c, x32, x33, x34, x35, x36_c, x38, x39, x40, x41_c, x42_c, x45_c, x46, x48, x50_c, x51_c, x54_c, x55, x56_c, x60_c, x61, x62, x63, x64_c, x65, x66, x67, x68_c, x70_c, x71, x72, x76, x77_c, x78_c, x79, x80, x81_c, x82, x83, x84_c, x85_c, x87_c, x88_c, x92, x93_c, x94, x95, x96, x98, x99);
and (w854, x0_c, x2_c, x4_c, x8, x11, x14_c, x17_c, x18_c, x19, x20_c, x22, x24_c, x25_c, x26, x27, x28, x32, x33, x35_c, x36, x39, x41_c, x45, x46, x47_c, x48_c, x49_c, x51_c, x52_c, x53, x54_c, x55, x56, x58_c, x59_c, x67_c, x68_c, x71_c, x73_c, x75_c, x76_c, x77, x78_c, x82_c, x83_c, x85, x87_c, x88_c, x89_c, x90, x93_c, x96, x97);
and (w855, x0_c, x3, x4_c, x5_c, x7, x8_c, x9_c, x10_c, x12, x17, x20, x22, x24, x26_c, x27_c, x28_c, x33, x38_c, x39_c, x42_c, x43, x44, x45_c, x46_c, x47_c, x48, x49_c, x51, x52, x54_c, x55_c, x57, x58_c, x59_c, x60_c, x61, x63_c, x64, x65, x70, x73_c, x74, x77_c, x78, x79, x80, x83_c, x85_c, x86, x88, x89_c, x93, x94_c, x95, x97_c, x98_c, x99);
and (w856, x0_c, x2_c, x4_c, x7_c, x9_c, x11, x12_c, x14_c, x15_c, x16_c, x17, x18_c, x19_c, x23, x25, x27, x28, x31, x33, x40_c, x41_c, x42, x44, x45_c, x48, x49_c, x50, x51, x52_c, x53, x56, x57, x58, x60_c, x61_c, x62, x67, x69_c, x70, x71, x74, x77_c, x78, x80_c, x82_c, x84_c, x86_c, x88_c, x90_c, x91, x92, x95_c, x97_c, x99);
and (w857, x9_c, x10_c, x16_c, x25_c, x44_c, x50, x57, x63_c, x64_c, x65, x68_c, x70, x83_c, x89, x92_c);
and (w858, x0_c, x1_c, x2_c, x3_c, x4_c, x6, x7_c, x8_c, x9, x11, x12, x17, x19_c, x20_c, x21, x22, x24_c, x25_c, x27_c, x29_c, x30_c, x31_c, x32, x33, x37_c, x39, x42, x44, x45, x46_c, x49, x50, x51_c, x52_c, x53_c, x55, x57, x61_c, x63, x66, x67_c, x69_c, x70, x72, x73_c, x76, x77_c, x79, x80_c, x81, x83_c, x85_c, x87, x88_c, x90_c, x92, x96, x98_c);
and (w859, x0, x1_c, x3_c, x7_c, x8_c, x9_c, x10, x11, x12, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x21_c, x22_c, x23_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29, x30_c, x31_c, x32, x33, x34, x35_c, x36, x37, x38_c, x39_c, x40, x41_c, x42_c, x43, x45, x47_c, x48, x49_c, x50, x51, x52, x53_c, x54_c, x55, x56_c, x57_c, x58_c, x59, x61_c, x63, x64, x65_c, x66, x67_c, x68, x69, x70, x71, x72, x73, x74, x75_c, x76_c, x77_c, x78_c, x79, x80_c, x81, x82_c, x83_c, x84, x85, x86, x88, x89, x90, x91, x92_c, x93_c, x94, x95, x96_c, x97, x98);
and (w860, x0, x1_c, x13, x22, x24, x25_c, x30, x43, x46_c, x48, x54_c, x60_c, x61_c, x65, x66, x67_c, x75_c, x81_c, x83, x87_c, x89, x98, x99_c);
and (w861, x1, x2, x3, x7, x8_c, x9_c, x10_c, x11, x13, x15, x16, x18_c, x21, x22_c, x23, x26_c, x27_c, x29_c, x31, x32_c, x34, x37, x38, x39_c, x40, x41_c, x42_c, x43, x45, x49_c, x50_c, x51, x53, x56, x57, x58_c, x61_c, x62_c, x63, x64_c, x68_c, x69, x70, x72, x75_c, x76, x77, x79, x81_c, x84, x87, x92_c, x95, x97, x98_c);
and (w862, x0, x1, x2_c, x3_c, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13_c, x14_c, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22, x23, x24, x25_c, x26_c, x27, x28_c, x29_c, x30_c, x31, x32, x33, x34_c, x35_c, x36, x37, x38_c, x39_c, x40_c, x42_c, x43_c, x44_c, x45_c, x48_c, x49_c, x51, x52_c, x54_c, x55, x56_c, x58, x59, x60, x61, x62_c, x63_c, x64_c, x65, x66, x67_c, x68_c, x69, x70, x71_c, x72_c, x73, x74, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x82_c, x84, x85_c, x86, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93, x94, x95_c, x96_c, x97, x98_c, x99);
and (w863, x0_c, x2, x3_c, x4, x5, x6_c, x8_c, x11, x13, x14_c, x15_c, x16_c, x17, x18_c, x20, x21_c, x22_c, x24_c, x25_c, x26, x28_c, x29_c, x30_c, x34, x35_c, x36_c, x38, x41_c, x42_c, x43, x44_c, x47_c, x48_c, x50, x51, x52_c, x53_c, x54, x56, x57_c, x60, x61_c, x62_c, x63, x67, x68_c, x69_c, x70_c, x72_c, x73_c, x74_c, x76, x78, x79_c, x80, x84, x85, x86_c, x89_c, x91_c, x92, x93_c, x94, x95, x96_c, x98_c, x99_c);
and (w864, x3, x5_c, x14, x38_c, x39_c, x42_c, x45_c, x51_c, x54, x64_c);
and (w865, x7, x9, x10_c, x12, x14_c, x18_c, x19_c, x22, x23, x24, x26, x27, x34, x40, x46_c, x48_c, x53, x55, x57_c, x62, x63_c, x65, x70_c, x71, x72, x73, x74_c, x79, x80, x84, x86, x87_c, x89, x90, x92, x98_c, x99);
and (w866, x3_c, x5, x6, x8, x16, x17_c, x21_c, x23_c, x26, x27, x34_c, x36, x38_c, x54, x57_c, x58_c, x61, x63, x66, x67, x69_c, x71_c, x73_c, x77, x79, x93_c, x95, x97_c, x98_c);
and (w867, x1, x2_c, x3_c, x4_c, x5_c, x6, x8_c, x11_c, x12, x13, x14_c, x15, x17_c, x20, x21, x22, x24_c, x26, x28, x29_c, x30_c, x31, x32, x33, x34_c, x35, x36_c, x38, x39_c, x40, x41_c, x42, x43_c, x44, x45, x47, x48, x49_c, x50, x51_c, x53_c, x54, x55, x56, x57, x58_c, x60_c, x61_c, x62_c, x63, x64_c, x66_c, x67, x68, x72_c, x73, x74, x75_c, x76_c, x77, x78, x79_c, x80, x82, x84, x85, x86_c, x87_c, x91_c, x92, x93_c, x94_c, x96, x97_c, x98, x99);
and (w868, x14_c, x22, x41_c, x42, x76, x79_c, x87, x95, x96, x98_c);
and (w869, x2, x3_c, x4_c, x5, x6, x7_c, x8, x11_c, x12_c, x15_c, x17_c, x18, x20_c, x21_c, x23, x24, x25, x26, x28_c, x29_c, x30_c, x31_c, x33, x34_c, x35_c, x39_c, x40_c, x41, x42, x43, x44, x46_c, x48_c, x50_c, x51, x52, x53_c, x54_c, x55_c, x56, x57, x58, x60_c, x61, x62, x63, x64, x65_c, x66_c, x67_c, x68, x69, x70, x71, x72_c, x73, x74_c, x75, x76, x77, x78, x79_c, x80_c, x82, x83_c, x84, x85_c, x86, x88, x89_c, x90, x91, x92_c, x94_c, x95, x96_c, x97, x98);
and (w870, x0, x1, x2_c, x4_c, x6_c, x7, x8_c, x12, x13, x15, x16_c, x21_c, x25_c, x27_c, x28, x30, x31, x33_c, x34_c, x35, x37, x38_c, x39, x40, x42, x43, x44_c, x47_c, x49_c, x52, x54_c, x55, x56, x58_c, x59, x61_c, x62_c, x64, x66, x67, x68, x69, x70_c, x74, x75, x76, x77, x80, x81, x84, x85_c, x86_c, x90, x91_c, x94, x95, x97, x98);
and (w871, x1_c, x2_c, x3, x4, x5_c, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x12, x13, x14_c, x15_c, x17, x18, x19, x20_c, x21_c, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32, x33, x34_c, x35, x36_c, x37, x38, x39, x40, x41, x42_c, x43, x44, x45, x46, x47, x48, x49_c, x50_c, x51, x52, x53_c, x54, x55_c, x56_c, x57_c, x58_c, x59_c, x60, x61, x62, x63, x64_c, x65, x66, x67, x68_c, x69, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78, x79_c, x80, x82, x83_c, x85_c, x86_c, x87_c, x88, x89, x90, x92_c, x93_c, x94, x95_c, x96, x97, x98);
and (w872, x0_c, x1_c, x2, x3_c, x4_c, x6, x7, x8, x9, x10_c, x12_c, x14_c, x15_c, x16, x17_c, x19_c, x20, x23, x24, x25, x27, x28_c, x29_c, x30_c, x31_c, x32, x33, x34, x35, x37_c, x38_c, x39, x40_c, x41, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x51, x52_c, x54, x56, x57, x58, x60, x61_c, x62, x63, x67, x69, x72_c, x73, x77, x78, x79_c, x80, x81_c, x83, x84_c, x85, x87_c, x88, x90, x92_c, x93, x94, x95, x97_c, x98_c);
and (w873, x1, x4_c, x5_c, x6, x7, x8, x10_c, x11_c, x12, x14_c, x15_c, x17_c, x18, x19_c, x22_c, x23, x24, x25, x26_c, x27_c, x28_c, x31, x32, x33, x36, x37_c, x38_c, x39_c, x40, x41_c, x43_c, x44_c, x45_c, x46_c, x47, x48_c, x49_c, x50, x52_c, x54, x55, x56, x57_c, x58, x59_c, x60, x61_c, x62_c, x63_c, x64, x66, x67, x68, x69, x72_c, x73_c, x74_c, x76, x78, x79_c, x81_c, x83_c, x84, x85, x86_c, x87, x88, x89, x90, x91_c, x93, x94, x95_c, x96_c, x97_c);
and (w874, x0, x2, x3_c, x9_c, x14, x15, x21, x25, x26_c, x28, x29_c, x31, x33_c, x35_c, x38, x41_c, x46, x55_c, x63_c, x65, x70_c, x91, x93_c, x95_c);
and (w875, x18, x42_c, x45, x51, x58);
and (w876, x1, x3_c, x4_c, x7_c, x9_c, x11, x19, x23_c, x27, x28, x29_c, x36, x37, x40, x42_c, x46_c, x48_c, x49, x50, x52, x55, x57, x58_c, x62_c, x64_c, x65, x67_c, x69, x70_c, x74, x76, x80_c, x85, x87_c, x90_c);
and (w877, x0_c, x1_c, x4, x6, x7, x8, x9_c, x10_c, x11_c, x15_c, x16, x18_c, x20, x21, x22_c, x23, x24, x25_c, x27, x28_c, x29, x30, x32, x34, x36_c, x37_c, x38_c, x39_c, x40_c, x41, x42, x43_c, x44, x46_c, x47, x48_c, x49, x50_c, x52_c, x54_c, x55_c, x56, x57, x59, x60, x62, x64, x65, x67, x68, x71_c, x72_c, x73, x74, x76, x77, x80, x81, x82, x83, x84, x87, x90_c, x91, x92, x93_c, x94, x95_c, x96, x97, x98, x99_c);
and (w878, x4, x5_c, x6_c, x7, x13, x18_c, x19, x20_c, x21_c, x22_c, x29_c, x33, x34, x35_c, x37, x38, x39_c, x42, x49, x50_c, x51_c, x52, x54, x58_c, x59, x60_c, x63, x66, x67, x70, x71_c, x73_c, x74, x75, x76, x77, x81, x83, x84, x85, x86_c, x93_c, x94_c, x96, x97);
and (w879, x0, x1_c, x2, x3, x4_c, x5_c, x6, x7, x11_c, x12, x13, x14_c, x15_c, x16, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36, x38, x39, x40_c, x41, x42, x43, x44_c, x45, x46_c, x47_c, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55_c, x56, x57_c, x58_c, x59_c, x60_c, x61, x62_c, x63, x64_c, x65_c, x66, x67_c, x68, x69_c, x70, x71, x72_c, x73_c, x74, x75, x76_c, x77_c, x78_c, x79, x80, x81, x82, x83, x84, x85, x86_c, x87_c, x88, x89_c, x90_c, x91, x92_c, x93_c, x94_c, x95, x96, x97, x99_c);
and (w880, x0_c, x1_c, x3, x4, x7, x9_c, x12_c, x13_c, x16, x26, x27_c, x30, x32, x34_c, x35_c, x39, x43, x45_c, x48, x49_c, x50_c, x52, x55_c, x58, x59, x66, x67, x71, x74_c, x77, x83, x85_c, x88_c, x89, x90_c, x92, x95_c, x97);
and (w881, x1_c, x3, x7, x8, x9_c, x10, x11_c, x13_c, x14_c, x15_c, x16, x17_c, x18, x20, x21_c, x24_c, x25, x28_c, x30, x36_c, x37, x41, x44_c, x48, x54, x58, x59, x62_c, x66_c, x68, x69, x71_c, x72, x73_c, x80_c, x82, x86_c, x87, x95);
and (w882, x0, x2, x3_c, x6_c, x8_c, x9, x10_c, x11, x13_c, x15, x16, x17, x18_c, x19_c, x20_c, x21, x24_c, x25_c, x26, x27_c, x28, x29, x30, x32, x33, x34, x35_c, x38_c, x40, x41, x44, x45, x46, x47, x48_c, x50, x51, x53_c, x55_c, x57_c, x59_c, x60_c, x61_c, x62_c, x63_c, x64, x68_c, x69, x70_c, x71_c, x72_c, x73, x74, x76_c, x77_c, x81, x82_c, x83, x84, x85, x87_c, x89_c, x90_c, x91_c, x93, x97, x99);
and (w883, x2_c, x4, x6, x7_c, x10_c, x11_c, x13, x17, x18, x30_c, x31, x38, x40_c, x41, x43, x48, x50, x52, x53_c, x55, x57, x63, x65_c, x68, x69, x72, x75, x77, x79, x84_c, x85, x89, x92, x94_c, x95_c, x97, x99_c);
and (w884, x3_c, x7_c, x12, x13_c, x14, x16, x18, x19_c, x23, x24_c, x25, x29, x34_c, x37, x38, x40, x43_c, x45, x48_c, x50_c, x52_c, x57, x59_c, x61_c, x64_c, x66, x68, x69_c, x74, x82, x84_c, x87_c, x89, x90_c, x92, x94_c, x97_c);
and (w885, x10_c, x35, x49_c, x64_c, x95_c);
and (w886, x1, x2, x3_c, x6_c, x9_c, x10, x11_c, x14_c, x17, x18_c, x20, x22_c, x24_c, x28, x29_c, x32_c, x36_c, x38, x39, x42_c, x45, x46_c, x47_c, x48_c, x49_c, x50_c, x52_c, x56, x59, x60_c, x61, x62_c, x65_c, x66_c, x67_c, x68, x73_c, x77, x78_c, x79_c, x85_c, x86, x87, x88, x91, x92, x93_c, x96, x97_c, x98, x99_c);
and (w887, x0_c, x2_c, x3, x5_c, x6, x7, x8, x9, x10, x11_c, x14, x15_c, x16, x17, x20, x21, x22, x23_c, x25, x26, x27, x28, x29, x30_c, x32, x33, x34, x36, x38_c, x40_c, x42_c, x43_c, x44, x46_c, x47, x48_c, x49_c, x50_c, x51_c, x52, x53, x54, x55, x60_c, x61, x62_c, x63_c, x64, x65, x67, x68_c, x72_c, x73, x74_c, x77, x78_c, x79, x80, x84_c, x85, x86, x88, x90_c, x92, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w888, x0_c, x3_c, x6, x11_c, x14, x15, x20, x22, x24, x25, x27_c, x29_c, x30_c, x33_c, x35, x39_c, x41_c, x44, x45_c, x46, x48_c, x51_c, x53, x55, x58_c, x60_c, x62_c, x63, x64, x65, x66_c, x67, x70_c, x72, x75_c, x85_c, x88, x89_c, x90, x91_c);
and (w889, x0, x1_c, x2, x3_c, x4_c, x5_c, x6, x7, x8_c, x10_c, x11, x12_c, x14_c, x15, x16, x17_c, x18, x19, x20_c, x21, x22_c, x23_c, x24_c, x25, x27, x28_c, x29, x30_c, x31_c, x32, x33_c, x34, x35_c, x36, x37, x40_c, x41, x42, x43_c, x44, x45, x46_c, x47, x48, x49_c, x50_c, x51, x52, x53_c, x54_c, x55, x56_c, x57_c, x58, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x69_c, x70, x71, x72_c, x73_c, x74_c, x76, x78, x79_c, x80, x81_c, x83, x84_c, x85_c, x86, x87, x88, x89_c, x90_c, x91_c, x92, x93_c, x94, x95, x96_c, x97, x98, x99_c);
and (w890, x0_c, x1_c, x2, x3, x4, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x14, x15_c, x16_c, x17_c, x19_c, x20, x21, x22_c, x23, x24_c, x25, x26, x27, x29, x30_c, x31, x32_c, x33, x34, x35_c, x36_c, x38, x39, x40_c, x41_c, x42, x43, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x54, x55_c, x57_c, x58, x59_c, x60_c, x61_c, x62, x63_c, x64_c, x65, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74, x76_c, x77, x78_c, x79_c, x80, x81, x82_c, x83_c, x84, x85_c, x86, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95_c, x97_c, x98, x99);
and (w891, x2, x10_c, x12_c, x17, x19, x29_c, x31_c, x34_c, x49_c, x50_c, x55_c, x59_c, x72_c, x73, x74, x75, x80, x82, x89_c, x97, x98_c);
and (w892, x0, x1_c, x2_c, x3, x4_c, x5_c, x6_c, x8, x9, x10, x11, x12, x13, x14_c, x15, x16, x17, x18_c, x19_c, x20, x21, x22_c, x23_c, x24_c, x25, x26_c, x27, x28_c, x29, x30_c, x31, x32_c, x33_c, x34, x35_c, x36, x37, x38_c, x39_c, x40, x41, x42, x43_c, x44, x45_c, x46_c, x47, x48, x49_c, x50_c, x51_c, x52, x53, x54, x55_c, x56_c, x57, x58, x59, x60, x61_c, x62_c, x63_c, x64, x65, x66, x67, x68_c, x69, x70_c, x71, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78, x79_c, x80, x81_c, x82_c, x83_c, x85, x86_c, x87_c, x88_c, x89_c, x90_c, x91, x92, x93, x94_c, x95, x96_c, x97, x98_c, x99_c);
and (w893, x0, x1, x2, x3, x4, x5, x6_c, x7_c, x8_c, x9_c, x10_c, x11, x12, x13_c, x14_c, x15_c, x16, x17_c, x18, x19_c, x20, x21, x22, x23, x24, x25_c, x26_c, x27, x28, x29_c, x30, x31, x32, x33_c, x34, x35, x36, x37_c, x38, x39, x40_c, x41_c, x42_c, x43, x44_c, x45, x46, x47, x48_c, x49, x50, x51, x52_c, x53, x54, x55, x56, x57, x58, x59_c, x60, x61_c, x62, x63_c, x64_c, x65_c, x66, x67, x68_c, x69_c, x70, x71_c, x73_c, x74_c, x75, x76_c, x77, x78_c, x79_c, x80_c, x81, x82, x83_c, x84, x85, x86_c, x87_c, x88_c, x89, x90, x91_c, x92, x93_c, x94, x95, x96, x97_c, x98, x99_c);
and (w894, x1, x3_c, x7, x12_c, x13, x14, x15_c, x20_c, x21_c, x22, x25_c, x26, x28, x33_c, x37, x46, x48_c, x50, x55, x62, x64, x65, x72, x75, x81, x84, x90_c, x93, x95_c);
and (w895, x1, x6, x7_c, x12_c, x13, x22_c, x23_c, x25_c, x27, x28_c, x31, x32_c, x33_c, x37_c, x39_c, x40_c, x43, x44, x49, x55_c, x58_c, x61, x63_c, x64_c, x67_c, x68, x70, x75, x78_c, x88, x89_c, x90, x91_c, x94, x98);
and (w896, x8_c, x11_c, x12_c, x14, x15_c, x19_c, x24, x26_c, x28_c, x32_c, x33_c, x39_c, x40, x47, x48_c, x57_c, x66, x69, x70, x76, x77_c, x91_c, x95_c, x98);
and (w897, x0_c, x1, x2_c, x3, x4_c, x6, x7, x8_c, x12_c, x13, x14_c, x15, x16, x17, x20, x21_c, x23_c, x24, x25, x26, x27_c, x28_c, x30_c, x31_c, x33, x34_c, x35_c, x36_c, x37_c, x38_c, x40, x42, x43_c, x44, x45_c, x46_c, x49_c, x50_c, x51_c, x52, x53, x54, x55_c, x57, x58_c, x63, x64, x65_c, x66_c, x67, x69, x71, x72_c, x73, x74, x75, x76_c, x77_c, x78_c, x79_c, x84_c, x88_c, x90, x91, x92, x93, x94_c, x95, x96_c, x98, x99_c);
and (w898, x2_c, x3, x6_c, x8, x11_c, x12, x16, x19_c, x27_c, x31, x33_c, x37, x43, x47_c, x50, x51, x60, x63_c, x64, x65_c, x67_c, x68_c, x69, x70_c, x71_c, x72, x75_c, x76, x78, x80, x81_c, x87_c, x90_c, x92, x95_c);
and (w899, x1, x2_c, x3_c, x8_c, x12, x13, x17_c, x18, x22_c, x23_c, x27_c, x29, x31_c, x35_c, x39, x40_c, x41, x44, x48, x52_c, x53, x55_c, x56, x58_c, x68_c, x73, x77, x78_c, x80, x84, x90_c, x93_c, x95_c, x96, x98, x99);
and (w900, x2, x6, x7, x12_c, x14_c, x29_c, x31, x32, x33_c, x34_c, x35, x36, x37_c, x40, x41_c, x43, x44, x45, x46_c, x47, x53_c, x55, x56_c, x65, x74, x75, x76_c, x78, x81_c, x82, x83_c, x86, x87, x88_c, x90, x91, x92_c, x95_c, x97);
and (w901, x1, x2_c, x7, x9_c, x10_c, x12, x13_c, x14, x15_c, x16_c, x18, x19, x21, x23_c, x27_c, x29_c, x31_c, x33_c, x34, x35, x38_c, x41_c, x42, x45, x46_c, x47_c, x48_c, x50, x52, x53_c, x56, x58_c, x59_c, x60, x62_c, x63, x64, x66_c, x69_c, x70_c, x71_c, x74, x75, x76, x78, x79_c, x86, x87_c, x88_c, x89, x90, x91_c, x92, x93, x94, x95, x96, x97);
and (w902, x5, x7_c, x15_c, x17, x31, x34, x38_c, x40, x41, x47, x67, x69_c, x70_c, x76, x79_c, x85_c, x87_c, x88_c, x91, x94);
and (w903, x0, x1, x2, x3_c, x4, x5, x6_c, x7_c, x8_c, x9, x10_c, x11, x12, x13, x14, x15_c, x16, x17, x18_c, x19_c, x20_c, x21_c, x22_c, x23, x24, x25_c, x26, x27_c, x28, x29, x30, x31, x32_c, x33, x34, x35_c, x36, x37, x38, x39, x40, x41_c, x42_c, x43, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56, x57, x58, x59_c, x60_c, x61_c, x62, x63_c, x64, x65_c, x66, x67, x68, x69, x70_c, x71_c, x72, x73, x74, x75, x76_c, x77_c, x78_c, x79, x80_c, x81, x82, x83, x84_c, x85_c, x86_c, x87, x88, x89_c, x90, x91, x92_c, x93, x94_c, x95, x96_c, x97_c, x98_c, x99);
and (w904, x11_c, x14_c, x16, x18_c, x24_c, x31_c, x38, x43_c, x45, x47_c, x48_c, x52_c, x62, x65, x70_c, x80, x83_c, x86_c, x87_c, x89_c, x95, x99_c);
and (w905, x0_c, x1, x2_c, x3, x4_c, x5, x6_c, x7_c, x8_c, x9_c, x10, x12_c, x15, x16, x17, x18, x19, x20, x21, x22, x23_c, x24_c, x25_c, x26_c, x28_c, x29, x30, x31, x32_c, x33_c, x34, x35_c, x36, x37_c, x38, x39_c, x40, x41_c, x42_c, x43_c, x44, x46_c, x50, x51, x52, x53, x54_c, x55, x56_c, x58_c, x59_c, x60_c, x61_c, x62_c, x63, x66_c, x67_c, x68, x69_c, x70, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78, x79, x80_c, x81, x82, x83_c, x84, x85, x87_c, x88, x89, x90, x91_c, x92_c, x93, x94, x95, x97_c, x98_c, x99_c);
and (w906, x12_c, x14, x20_c, x26, x44, x53_c, x74, x99);
and (w907, x2, x3, x4, x6_c, x7_c, x8, x9, x10, x12_c, x16, x17_c, x18_c, x20_c, x21, x22_c, x24_c, x25, x27_c, x28_c, x29_c, x30_c, x32, x34_c, x35_c, x36, x38_c, x40_c, x41, x44_c, x45, x46, x47_c, x50, x51_c, x52_c, x55_c, x56_c, x57, x58, x60, x61_c, x65_c, x66, x67_c, x68_c, x69_c, x70_c, x72, x75, x76, x77_c, x78_c, x79, x80, x81, x82_c, x85_c, x86_c, x87, x88_c, x89, x91, x92_c, x94_c, x95_c, x96, x97_c, x98_c);
and (w908, x0, x1, x3_c, x4, x5_c, x8, x9_c, x11, x13, x15, x17_c, x18_c, x20_c, x21_c, x22_c, x23_c, x24_c, x25_c, x26, x27, x28, x29, x30, x32, x35_c, x36, x37_c, x38_c, x39, x41, x42, x43, x44, x45_c, x47_c, x49_c, x50, x51, x52, x53, x54_c, x55_c, x57, x59, x60, x61, x62_c, x63_c, x64_c, x65_c, x66, x68_c, x69_c, x71_c, x72, x73, x74, x75, x76_c, x77, x78, x79_c, x80, x81, x84, x85_c, x86, x87, x89_c, x90, x91, x92_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w909, x2_c, x4, x6, x9_c, x10, x18_c, x29, x30_c, x32_c, x38, x39_c, x40, x44, x52, x53_c, x54, x55, x57_c, x61_c, x62_c, x66, x70_c, x73, x75_c, x76_c, x87_c, x88_c, x91, x99);
and (w910, x0, x1, x2, x3, x4, x5, x6_c, x7_c, x8_c, x9, x10, x11, x12, x13, x14_c, x15, x16_c, x17, x18, x19, x20_c, x21, x22, x23, x24_c, x25_c, x26, x27_c, x28, x29_c, x30_c, x31, x32_c, x33_c, x34, x35_c, x36_c, x37_c, x38, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x47, x48, x49, x50, x51_c, x52, x53_c, x54, x55_c, x57, x58, x59_c, x60, x61, x62_c, x63, x64, x65, x66_c, x67, x68, x69, x70_c, x71, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x81_c, x82_c, x83, x84_c, x85_c, x86, x87_c, x88, x89_c, x90, x91_c, x92, x93_c, x94_c, x95, x96, x97_c, x98, x99);
and (w911, x0, x1, x2_c, x3_c, x4_c, x5_c, x6_c, x7_c, x11, x12, x13_c, x15_c, x17, x18, x20_c, x21_c, x22_c, x23_c, x24_c, x25, x28_c, x29_c, x31_c, x32, x33_c, x34_c, x35, x36_c, x37, x38, x39, x40_c, x42, x43_c, x44, x45_c, x46_c, x47, x48_c, x49_c, x50, x51, x52_c, x53, x54, x55, x56, x58_c, x59, x61_c, x62, x64_c, x66, x67_c, x68, x69, x70, x72, x73_c, x75_c, x76, x80, x81_c, x82_c, x84_c, x85, x88_c, x89_c, x91_c, x94_c, x95, x96, x97);
and (w912, x10_c, x27_c, x31, x35_c, x37, x62_c, x63_c, x65, x67, x68, x69, x73, x74_c, x85, x89, x95_c, x98_c);
and (w913, x3_c, x4, x8, x10, x14_c, x16, x19_c, x24, x29, x33, x34, x35_c, x38, x42, x43_c, x47_c, x48, x49, x50, x52_c, x53_c, x58, x60, x61_c, x63, x64, x65, x71_c, x74_c, x76_c, x77_c, x80_c, x81, x82, x87, x90, x92_c, x95, x96);
and (w914, x2_c, x3_c, x4_c, x5, x7, x8_c, x9_c, x10, x11_c, x13_c, x14_c, x15_c, x16_c, x17, x18, x19_c, x21_c, x22, x24, x26_c, x28_c, x29, x30, x31_c, x32_c, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40, x42, x43, x44_c, x45, x46_c, x47, x49_c, x50_c, x51_c, x52, x53_c, x55_c, x56_c, x57_c, x58, x59_c, x60_c, x64, x65, x66, x67_c, x68, x70, x72_c, x73_c, x74, x75_c, x76_c, x77_c, x78, x79, x80_c, x81_c, x82, x84, x86_c, x87, x88_c, x90_c, x91, x94_c, x96, x97, x98);
and (w915, x1, x2_c, x3, x4, x5, x8_c, x9, x11_c, x12, x13, x15_c, x17, x18, x19, x21, x22_c, x23_c, x25, x29_c, x34, x37, x38_c, x39_c, x40, x41_c, x43_c, x45, x46_c, x49_c, x52, x53, x55_c, x56_c, x57, x58, x60, x61_c, x64_c, x69, x72, x74_c, x76, x77, x79, x80_c, x84, x86, x87, x88, x89, x91, x92, x93, x94, x96, x97, x98, x99_c);
and (w916, x0, x1, x2, x3_c, x4_c, x5, x6, x9_c, x10_c, x12_c, x13_c, x14_c, x15_c, x17, x19, x20, x21, x22, x23_c, x24_c, x26, x27_c, x29, x30, x31_c, x33, x34, x36_c, x37_c, x40_c, x43_c, x45_c, x46_c, x47_c, x49, x50_c, x54_c, x55_c, x56, x57, x59_c, x60_c, x61_c, x62, x64, x65, x67, x69_c, x70, x73_c, x74_c, x75_c, x78, x79_c, x80, x81_c, x82_c, x83, x84, x86_c, x87, x88_c, x89_c, x92, x93, x95_c, x96_c, x97);
and (w917, x1, x3, x4_c, x5, x7, x8, x9, x10_c, x11_c, x14, x15, x16, x17, x18, x19, x23, x24, x26, x27_c, x28, x30_c, x31, x32, x34, x35_c, x36_c, x37, x40_c, x42_c, x43, x44_c, x47, x48_c, x49, x51_c, x52_c, x53_c, x54_c, x55, x57, x58_c, x59_c, x60, x61, x63_c, x65_c, x68, x71_c, x72_c, x75_c, x77_c, x78_c, x79_c, x81_c, x82, x84_c, x85, x86, x87, x88, x90, x91, x92_c, x94, x96, x99_c);
and (w918, x0_c, x1_c, x2, x3, x4_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12_c, x13, x14_c, x15, x16, x17_c, x18_c, x19, x20_c, x21_c, x22_c, x23_c, x24, x25, x26_c, x27_c, x28_c, x29, x30_c, x31, x32, x33, x34_c, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x43, x44, x45, x46, x47_c, x48_c, x49_c, x50_c, x51_c, x52_c, x53, x54_c, x55_c, x56_c, x57, x58_c, x59_c, x60, x61, x62_c, x63, x64, x65, x67, x68_c, x69, x70, x71, x72, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80_c, x81, x82, x83, x84_c, x85, x86_c, x87, x88, x89, x90, x91, x92_c, x93, x94_c, x95_c, x96_c, x97, x98_c);
and (w919, x0_c, x1, x2_c, x3_c, x4_c, x5, x6_c, x7_c, x8, x9, x10_c, x12, x13_c, x15_c, x17_c, x19, x20, x21_c, x22, x23_c, x24, x25, x26, x27, x28_c, x29_c, x30_c, x31, x32_c, x33_c, x34, x35, x36_c, x37, x38, x39_c, x40, x42_c, x43_c, x44_c, x45_c, x46, x47, x48_c, x49_c, x50, x51_c, x52, x53, x54, x55, x56_c, x57, x58, x59, x61, x62_c, x63_c, x64, x65_c, x66_c, x67, x68_c, x69_c, x70, x71_c, x72_c, x73_c, x74, x75_c, x76_c, x77, x78_c, x79_c, x80_c, x81, x83, x84, x85_c, x86_c, x87, x88, x89_c, x90_c, x91_c, x92_c, x94_c, x95_c, x96, x97_c, x98, x99_c);
and (w920, x8, x9_c, x11_c, x13, x16_c, x17, x18_c, x19, x23, x24, x25, x28_c, x30, x31_c, x33_c, x38, x39, x42, x43, x44, x45, x50, x51_c, x54, x56_c, x59, x63, x68, x69, x72_c, x74_c, x76_c, x79_c, x80_c, x81_c, x84_c, x86_c, x87, x89, x92, x94, x95, x97, x98);
and (w921, x5_c, x9, x12_c, x13, x14, x25_c, x32_c, x35_c, x47, x48, x50, x58_c, x63_c, x67_c, x75, x80, x86_c, x93, x94, x95_c, x96);
and (w922, x1, x2, x4, x9, x11, x12, x17, x21, x22_c, x23, x24, x26, x34, x35_c, x36, x37_c, x38_c, x39, x40, x41_c, x43_c, x44, x46_c, x49, x51, x54_c, x65, x66_c, x68_c, x72_c, x80, x85, x91_c, x93_c, x94, x95, x96_c, x98);
and (w923, x2_c, x52_c, x70_c);
and (w924, x0, x1, x3_c, x4_c, x5_c, x6_c, x7, x9_c, x10, x11, x14, x15, x16, x17, x18_c, x19, x20_c, x22_c, x23, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31_c, x32, x33_c, x34, x35, x36_c, x37_c, x38_c, x39_c, x41, x42_c, x43, x44, x45, x46_c, x47_c, x48, x49, x50_c, x52_c, x53, x54_c, x56_c, x58_c, x59, x60_c, x61, x62_c, x63, x64_c, x65, x66_c, x67, x68_c, x70, x71_c, x73, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80_c, x81_c, x82_c, x83, x84, x85, x86, x87_c, x88, x89, x90, x91_c, x92, x93, x94_c, x95_c, x96_c, x97, x98_c, x99_c);
and (w925, x0_c, x1_c, x3, x4_c, x5, x7_c, x8_c, x10, x11_c, x13, x14, x16, x18, x19_c, x22, x23_c, x24_c, x25, x26, x27_c, x28_c, x29, x30_c, x32, x33, x34_c, x35, x36, x37_c, x38, x39, x40_c, x41, x42, x43, x45, x46, x47, x49, x51_c, x53_c, x55, x56, x57, x58, x59, x63_c, x67, x68_c, x69, x70_c, x71, x72_c, x73, x75_c, x76, x77_c, x78_c, x80, x81, x82, x83_c, x84, x85_c, x86, x87_c, x89_c, x90, x93_c, x94, x96, x97, x99);
and (w926, x0, x1, x2_c, x6_c, x7_c, x8_c, x10, x12, x14_c, x15_c, x16_c, x17_c, x19, x20_c, x22, x24, x25_c, x27, x31_c, x32_c, x33, x34_c, x37_c, x38, x39_c, x40_c, x41, x42, x43, x44, x45, x46_c, x47_c, x48_c, x49_c, x50, x51_c, x53, x54, x55, x56_c, x57, x58, x60_c, x61, x62_c, x64_c, x66, x67_c, x70_c, x71_c, x72, x73, x75_c, x76_c, x80_c, x81_c, x83_c, x85_c, x92, x93_c, x99_c);
and (w927, x0_c, x2_c, x4, x5, x7_c, x9_c, x13_c, x14, x16_c, x18, x21, x23_c, x24_c, x25_c, x26, x27_c, x31, x34, x35, x37, x44, x45, x49, x50_c, x51, x52_c, x54, x59_c, x60, x61_c, x64, x65, x68, x70, x71, x73_c, x74, x78_c, x80_c, x81_c, x82, x86, x88, x92_c, x93_c, x94_c, x95_c, x97, x99_c);
and (w928, x0, x1_c, x2_c, x3_c, x4_c, x5, x6, x7_c, x8_c, x9_c, x10, x11_c, x12_c, x13, x14_c, x15, x16, x17_c, x18_c, x19_c, x20, x21, x22_c, x23, x24_c, x25_c, x26, x27_c, x28_c, x29_c, x30, x31, x32, x33_c, x34, x35_c, x36, x37_c, x38_c, x40, x41_c, x42, x43, x44, x45_c, x46_c, x47, x48, x50_c, x51_c, x52, x53, x54_c, x55_c, x56_c, x57_c, x58_c, x59, x60, x61, x62, x63, x64, x65, x66_c, x67_c, x68_c, x69, x70, x71, x72, x73, x74_c, x75, x76_c, x77, x78, x79, x81, x82, x83, x84_c, x85, x86_c, x87, x88_c, x89_c, x90, x91_c, x92_c, x93_c, x94_c, x95_c, x96_c, x97_c, x98, x99_c);
and (w929, x0, x2_c, x3_c, x5, x7_c, x9, x10_c, x11, x12, x13_c, x15, x18, x20_c, x23_c, x25, x26, x28, x31, x33_c, x37, x39, x40_c, x42, x47, x48, x49, x51, x52_c, x53, x54_c, x55_c, x57_c, x60, x62_c, x64, x67, x75, x76_c, x78, x80, x81_c, x82, x84_c, x86, x87_c, x88, x90, x95_c, x97, x98);
assign w930 = x83_c;
and (w931, x0, x1, x2_c, x3, x5_c, x7, x9, x10, x11_c, x13_c, x17, x18, x19_c, x20_c, x21, x25_c, x27, x28_c, x29, x32, x33_c, x35_c, x36, x42_c, x43_c, x44, x46, x48_c, x49_c, x51_c, x52_c, x54_c, x56, x58_c, x60, x63_c, x64, x66_c, x68, x70_c, x74, x75, x77_c, x80_c, x81_c, x82, x83, x86, x88, x89, x91_c, x92, x95, x97);
and (w932, x0, x1_c, x2, x3, x5, x8, x10_c, x11, x12_c, x13, x14, x15, x16, x17, x18_c, x20, x22, x24, x25_c, x27_c, x28_c, x29, x32, x33, x35_c, x38, x40_c, x41, x42_c, x43, x44_c, x47_c, x49, x51_c, x53_c, x54, x56, x58, x59_c, x60, x61_c, x62_c, x63, x64, x69_c, x70, x71, x73_c, x74, x75_c, x77, x78_c, x80, x81, x82_c, x83, x84, x85_c, x86, x87_c, x88, x89_c, x90_c, x94, x97_c, x98, x99);
and (w933, x26_c, x29_c, x31, x36_c, x38_c, x39, x47, x56, x63_c, x68_c, x78, x84_c, x86, x88_c, x89_c, x92, x93, x97);
and (w934, x0_c, x1_c, x2, x4, x5_c, x6, x7, x8_c, x9_c, x10, x11_c, x12_c, x13_c, x14_c, x15_c, x16_c, x17, x19, x20, x21, x22, x24, x27_c, x28, x29_c, x30_c, x31, x32, x33, x35_c, x36_c, x37, x38_c, x39, x40_c, x41, x44_c, x46_c, x47, x48_c, x49_c, x51, x53_c, x54_c, x55, x56_c, x60, x61_c, x62, x63_c, x66_c, x67, x68, x69_c, x70, x71_c, x72, x73, x75, x76, x77_c, x78_c, x79, x80, x81, x82, x83_c, x84, x85_c, x86, x87, x88_c, x89_c, x92, x93_c, x94_c, x95, x96, x97_c, x98_c);
and (w935, x0, x1_c, x2_c, x3_c, x4_c, x6_c, x8, x9_c, x10, x11_c, x12_c, x13_c, x14, x15_c, x16, x17_c, x20_c, x21_c, x22, x23, x24, x25, x27, x28_c, x29_c, x30_c, x31_c, x32_c, x33, x34, x35_c, x36, x37_c, x38_c, x39_c, x40_c, x41_c, x43_c, x44, x45_c, x48, x49_c, x50, x51_c, x53_c, x54, x55_c, x56, x58_c, x59, x60, x61, x62_c, x63, x64, x65_c, x66_c, x67_c, x68_c, x69, x70_c, x71, x73_c, x74, x75, x76_c, x78, x79_c, x80, x81, x82_c, x85, x86_c, x87_c, x88, x89_c, x90_c, x91, x93, x94, x95_c, x96_c, x97_c, x98_c, x99);
and (w936, x3, x4, x5_c, x6_c, x13_c, x14, x15, x17, x18_c, x20_c, x21, x23_c, x24_c, x25_c, x26_c, x29_c, x32, x35_c, x36_c, x37_c, x39, x41, x45, x46_c, x48_c, x49, x51, x52_c, x53_c, x55_c, x56_c, x57, x59, x62, x63, x64, x65_c, x67, x71, x72_c, x74_c, x76_c, x77_c, x78_c, x79_c, x81_c, x83, x84_c, x85_c, x89_c, x90_c, x92_c, x94, x95, x96_c, x98, x99);
and (w937, x1_c, x6, x8, x10, x20, x24, x27_c, x28, x29, x34, x35, x40, x43_c, x44, x45_c, x46_c, x48_c, x49_c, x53, x59_c, x61, x63, x67_c, x69_c, x70, x71_c, x77, x79_c, x80, x91, x96_c);
and (w938, x0, x1, x3, x4_c, x5_c, x6, x8_c, x10_c, x12_c, x13, x15, x16, x20_c, x21, x23, x27_c, x28_c, x29_c, x30_c, x32_c, x33_c, x34_c, x36_c, x37_c, x44_c, x45, x47_c, x48_c, x49_c, x52, x53, x55_c, x56_c, x57, x58, x59, x61, x63_c, x65, x68, x69, x70, x71_c, x72, x73, x76, x79_c, x80, x81_c, x82, x84, x87_c, x89, x93_c, x96, x97_c, x98);
and (w939, x0_c, x1_c, x2, x3, x4, x5, x6_c, x7, x8, x9_c, x10, x11_c, x12, x13, x14_c, x15_c, x17_c, x18, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x30_c, x31_c, x32, x33_c, x34_c, x35, x36, x37_c, x38, x39, x40, x42, x43, x44_c, x45, x46, x47_c, x48_c, x49, x50_c, x52, x53, x54, x55_c, x56_c, x57_c, x58, x59, x60, x62_c, x63, x64_c, x65, x66, x67, x69_c, x70_c, x71_c, x72, x73_c, x74, x75, x76_c, x77_c, x78_c, x79_c, x80_c, x82_c, x83, x84, x85_c, x86_c, x87, x88, x89_c, x91, x92, x93_c, x95_c, x96_c, x97, x98, x99);
and (w940, x1_c, x4, x5_c, x9, x13, x15_c, x18_c, x19, x21, x22_c, x26_c, x27, x30_c, x31_c, x32_c, x35, x38_c, x40, x46, x48_c, x49, x50, x51_c, x52, x55, x56, x57_c, x60_c, x72, x73, x76, x79, x82_c, x84, x85_c, x87, x88_c, x90_c, x91_c, x94_c, x98_c);
and (w941, x0, x1_c, x2_c, x3_c, x4, x7_c, x10, x11_c, x12, x13, x14_c, x15, x16_c, x18_c, x20_c, x21_c, x22_c, x23, x24, x25_c, x26_c, x27, x28_c, x29, x30, x31_c, x32, x33, x34, x35, x36, x37_c, x38_c, x39_c, x40, x41, x42_c, x43_c, x45, x46, x47, x48, x49_c, x50, x51_c, x52, x53_c, x54, x55, x56, x57, x58_c, x59_c, x60, x61_c, x62, x63, x65, x66_c, x67_c, x68_c, x69, x71, x72_c, x73, x75, x76, x77, x78, x79, x80, x81_c, x82_c, x83, x84_c, x85_c, x86, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94, x95, x96_c, x97_c, x98, x99);
and (w942, x0_c, x2_c, x3, x5_c, x9, x10, x11_c, x12_c, x15, x16_c, x17, x18_c, x19, x20, x21, x22_c, x23, x24, x25_c, x26_c, x28_c, x30, x31, x32_c, x33_c, x35_c, x36_c, x37_c, x39_c, x42_c, x43, x45_c, x49_c, x51, x53, x57, x60_c, x61_c, x63_c, x65_c, x66_c, x67, x68_c, x69, x71_c, x74, x76, x77_c, x79_c, x80, x82, x84_c, x85_c, x87, x93);
and (w943, x2, x4, x5_c, x6, x8_c, x10_c, x13, x16_c, x17_c, x21_c, x22_c, x23, x27, x34_c, x36_c, x38, x41_c, x42_c, x52_c, x56_c, x58, x59, x60, x61_c, x64, x65, x66, x68_c, x69_c, x71, x73, x75_c, x78_c, x83_c, x85, x86_c, x89, x90, x91, x92_c, x97_c, x98);
and (w944, x0, x1_c, x2, x4_c, x5_c, x6, x7, x8, x9, x11, x12, x13_c, x14, x16, x17, x18, x19_c, x21, x22_c, x23_c, x24_c, x25, x26, x27_c, x28_c, x29, x30_c, x31_c, x32, x34_c, x35_c, x36_c, x37_c, x38_c, x39, x40, x41_c, x43, x44, x45, x47_c, x48_c, x49, x50_c, x51_c, x52, x54, x56, x57, x58_c, x59_c, x60, x61, x62, x63_c, x64_c, x65, x66, x67, x68, x69, x70, x73_c, x74, x75, x76_c, x77_c, x78, x79_c, x80, x81_c, x82, x84_c, x85, x86_c, x87, x88_c, x90, x91, x92_c, x93, x94_c, x95, x96_c, x97_c, x98, x99_c);
and (w945, x3, x14, x21, x23_c, x24_c, x32_c, x33, x37_c, x38, x45, x59, x61, x70_c, x76_c, x77, x84_c, x87_c, x89, x92);
and (w946, x0_c, x2, x5, x6_c, x9, x11, x12_c, x14, x15, x18, x22, x25, x27_c, x32_c, x35_c, x36, x37, x39, x42, x45_c, x46, x47, x48_c, x50_c, x52, x53, x60_c, x64_c, x67, x68, x70, x71, x75_c, x76, x77_c, x79, x84_c, x87, x91, x98, x99);
and (w947, x4_c, x5, x6_c, x22, x31, x51_c, x59_c, x61, x64, x66, x70_c, x75_c, x79_c, x81_c, x82_c);
and (w948, x0_c, x1_c, x4_c, x5_c, x6, x8_c, x9, x10, x12_c, x13, x14, x16_c, x17_c, x18_c, x19_c, x20_c, x21, x22_c, x23_c, x24, x26, x27, x30_c, x31_c, x33, x36, x38, x41, x42_c, x44_c, x46_c, x50_c, x51_c, x54, x55_c, x56_c, x58_c, x59_c, x60_c, x61_c, x62, x63, x64_c, x67, x68, x70, x71, x72_c, x73, x74_c, x75, x78_c, x79_c, x80, x81_c, x82, x83_c, x87, x88_c, x89, x91_c, x94, x95_c, x96_c, x97);
and (w949, x0, x1_c, x2_c, x3_c, x4, x5, x6, x7_c, x8_c, x9, x10_c, x11, x12_c, x13, x15, x16, x17, x18_c, x19, x20_c, x21, x22, x23_c, x24_c, x25_c, x26_c, x27_c, x28, x29_c, x30_c, x31_c, x32, x33, x34, x35_c, x36_c, x37, x38_c, x39_c, x41, x42_c, x43_c, x44_c, x45, x46, x47, x48_c, x49, x50_c, x51, x52, x53_c, x54, x55, x56_c, x57_c, x59_c, x60, x61_c, x62_c, x63_c, x64_c, x65_c, x66, x67_c, x68_c, x69, x70_c, x71, x72, x73_c, x74_c, x75_c, x76, x77_c, x78, x79_c, x80, x81_c, x82, x83_c, x84, x85_c, x86_c, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94_c, x95, x96, x97, x98, x99);
and (w950, x0, x1, x3, x4_c, x5, x6, x7, x8_c, x9_c, x11_c, x12_c, x13, x14, x15, x18_c, x19_c, x20_c, x22, x23, x24, x25, x27, x28, x29_c, x30, x31, x32_c, x33_c, x34, x35_c, x38_c, x39, x40, x41, x42_c, x43_c, x44_c, x45, x46_c, x47_c, x48_c, x49, x50_c, x51, x52, x53_c, x55_c, x56_c, x57, x58_c, x59_c, x60, x61_c, x62_c, x63, x65_c, x66, x67_c, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x79, x80, x81, x82, x83, x84_c, x85_c, x86_c, x87_c, x88, x89, x90, x91, x92_c, x94_c, x95, x96_c, x97, x99_c);
and (w951, x0_c, x1, x3_c, x4_c, x5, x6_c, x7_c, x10_c, x11, x12_c, x13, x14_c, x15_c, x16, x17_c, x18_c, x19, x21_c, x23_c, x24, x27, x28_c, x29, x30, x32_c, x34_c, x35, x36_c, x37, x38, x39, x40, x41_c, x42, x43_c, x44, x45, x46, x47_c, x48, x50, x51, x52, x54, x55, x56, x57_c, x58_c, x59_c, x60_c, x61, x62, x63_c, x65, x66, x67_c, x69_c, x70, x71_c, x72_c, x73_c, x75, x76_c, x78, x80_c, x81, x82, x83, x84, x85, x86, x87_c, x88, x89_c, x90_c, x91, x92_c, x93, x94, x95_c, x96, x97_c, x99);
and (w952, x1, x4, x5, x8_c, x14_c, x16_c, x17, x19, x20_c, x23_c, x24_c, x25_c, x27_c, x30_c, x31_c, x35, x36_c, x37_c, x40, x43, x47_c, x48, x51, x54_c, x57, x58, x59_c, x60, x62_c, x66_c, x67, x70_c, x72_c, x79_c, x84, x92_c, x94, x95, x96, x97, x98_c, x99_c);
and (w953, x7_c, x26, x35_c, x40, x46_c, x53, x62, x66_c, x68_c, x71, x88_c, x92_c);
and (w954, x5_c, x9, x10, x11, x18_c, x26_c, x27_c, x32_c, x35_c, x38_c, x48_c, x50_c, x56, x61, x62_c, x67_c, x68_c, x74_c, x76, x80_c, x82, x84, x93_c);
and (w955, x2_c, x3_c, x4, x6, x9, x11_c, x12, x13, x14_c, x15, x16_c, x18, x19_c, x20_c, x22_c, x24_c, x25_c, x26_c, x27_c, x28_c, x29_c, x31, x32, x34, x35, x36_c, x37, x38_c, x39_c, x41_c, x43, x45, x46_c, x49, x50_c, x51_c, x52_c, x54, x55, x56_c, x58, x60_c, x62_c, x63_c, x64, x66_c, x67_c, x69_c, x70, x71_c, x74, x76_c, x77_c, x78, x81, x82_c, x83, x84_c, x85_c, x86, x87_c, x89, x90, x91, x92, x93, x94_c, x95_c, x96, x97_c, x99);
and (w956, x0, x7, x8_c, x10, x15_c, x26, x35, x36_c, x38, x40_c, x41, x43, x52, x59_c, x61, x63_c, x65_c, x66, x68_c, x70, x71, x73, x76, x78_c, x84, x85, x88_c, x93, x99);
and (w957, x2_c, x9, x12_c, x14, x17_c, x20, x23_c, x28_c, x41_c, x46, x53_c, x63, x64_c, x75, x79_c, x80_c, x82_c, x84, x92, x93_c);
and (w958, x0_c, x1_c, x2, x3_c, x5_c, x6, x7, x9_c, x10, x11_c, x12_c, x13_c, x15, x16, x17_c, x18_c, x19_c, x20, x21_c, x22, x23_c, x24_c, x25_c, x26_c, x27, x28, x29, x30_c, x31, x32, x33, x34_c, x35_c, x36_c, x37, x39_c, x40, x41, x42_c, x43_c, x44, x45_c, x46_c, x47_c, x48_c, x49, x50, x51_c, x52, x54_c, x55_c, x56, x57, x58_c, x59, x60, x62_c, x63_c, x64_c, x65_c, x66_c, x67_c, x68_c, x69_c, x70_c, x71_c, x72, x73, x74, x75, x76, x77_c, x78, x79_c, x81_c, x83_c, x85_c, x86_c, x87_c, x88_c, x89, x90_c, x91_c, x92_c, x93_c, x94_c, x95, x96, x97_c, x98, x99_c);
and (w959, x0, x7_c, x9, x12, x21_c, x34, x36_c, x39_c, x44_c, x49, x50, x52_c, x60_c, x66, x75, x76_c, x80, x81_c, x82_c, x86, x92_c, x93);
and (w960, x3_c, x4, x6, x8, x10, x11_c, x12_c, x14_c, x17, x20_c, x21_c, x22_c, x23, x25, x26_c, x27, x30, x31_c, x32, x33, x35_c, x36, x38_c, x40_c, x41, x42, x48, x49, x50, x51_c, x53_c, x58, x59_c, x60, x62, x64, x66_c, x68, x69_c, x71, x73, x74, x76, x78_c, x79, x80_c, x81_c, x82_c, x83_c, x84_c, x85_c, x87, x88_c, x89, x90_c, x91, x92, x93, x96, x99_c);
and (w961, x3_c, x4_c, x6, x9_c, x10_c, x12_c, x13_c, x19, x20_c, x21_c, x24, x28, x31_c, x32_c, x33_c, x39, x40, x41_c, x42, x45, x47, x56, x57, x60, x62, x63, x69_c, x70, x72, x75_c, x76, x79_c, x81_c, x83, x84, x91_c, x95_c, x96_c, x97);
and (w962, x2_c, x3_c, x4_c, x6_c, x9, x10_c, x12_c, x13, x14, x15_c, x17_c, x18_c, x19_c, x21_c, x24_c, x25, x26, x27, x29_c, x30, x32_c, x33, x35, x36, x37_c, x39, x40_c, x45_c, x48_c, x50_c, x52_c, x56, x58, x59, x60_c, x61, x65_c, x67_c, x68_c, x69_c, x70, x71, x72, x73, x77_c, x78_c, x79, x81_c, x83_c, x85, x88_c, x89, x90, x91_c, x92_c, x93, x95_c, x97_c);
and (w963, x0, x1_c, x4_c, x9, x10_c, x12_c, x13_c, x15_c, x16_c, x19_c, x20, x21, x22, x23, x28, x29_c, x31_c, x32_c, x34_c, x35_c, x37_c, x38, x44, x47, x50, x53_c, x55, x56, x57, x61, x62_c, x64, x65_c, x66_c, x69, x70, x74_c, x77_c, x78, x80_c, x82, x85, x87, x90_c, x93, x94_c, x96_c, x97_c, x98);
and (w964, x0_c, x4_c, x11, x14_c, x16, x17, x24_c, x25_c, x28, x29, x36_c, x37_c, x39_c, x51, x53, x55, x58, x59, x61, x69_c, x71_c, x74_c, x75, x76_c, x78_c, x79_c, x81, x82_c, x84, x87, x88, x95_c, x97_c, x98_c, x99);
and (w965, x3_c, x5, x6_c, x9, x10_c, x14_c, x15_c, x24, x25, x27, x29_c, x31, x32_c, x34, x35_c, x37, x38, x41, x43, x44_c, x46, x48, x50, x51, x53_c, x54, x57_c, x58_c, x62, x63_c, x68_c, x69_c, x71_c, x72, x73, x77, x78_c, x79_c, x80, x82_c, x83_c, x84_c, x85, x86_c, x88_c, x90_c, x92, x93);
and (w966, x0, x2, x3, x5, x7_c, x8, x10_c, x12_c, x13_c, x15, x17_c, x18, x19, x20, x22, x23_c, x24, x25, x26, x27_c, x28, x29, x31_c, x32_c, x35, x36, x39_c, x40, x41, x42_c, x43_c, x44, x45, x46_c, x48_c, x49_c, x51_c, x52, x53_c, x54, x55, x56, x58, x59, x60_c, x62, x63_c, x64, x65_c, x66, x67_c, x68, x69_c, x72_c, x73_c, x74_c, x75, x76_c, x77_c, x78, x79, x80_c, x81, x82_c, x83, x84, x85, x86, x87, x88_c, x89_c, x90, x91, x92, x93, x94, x95_c, x97, x98_c, x99);
and (w967, x0_c, x1_c, x3_c, x5_c, x6_c, x7_c, x9_c, x10, x12, x13, x14_c, x15_c, x16, x17, x18_c, x20_c, x21, x23_c, x24, x25_c, x29, x31, x32, x33_c, x34, x35_c, x36_c, x38, x41_c, x42, x44_c, x45, x47_c, x48_c, x49_c, x50, x51_c, x52_c, x54_c, x55_c, x56_c, x60, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x70_c, x72_c, x73, x74_c, x75_c, x76, x77_c, x78, x79, x81_c, x82_c, x84, x85_c, x87_c, x88, x89, x90_c, x92_c, x93_c, x94_c, x95_c, x97, x98_c);
and (w968, x0, x1, x2, x3, x4, x5_c, x6_c, x7, x8_c, x9, x10_c, x11, x12, x13_c, x14_c, x15_c, x17_c, x24, x25, x26_c, x29_c, x30_c, x31, x32_c, x33, x34_c, x35, x36, x37, x38_c, x41, x42_c, x43, x44_c, x46_c, x47_c, x48_c, x49_c, x50_c, x53, x54_c, x55, x57_c, x58, x59_c, x61, x62, x63_c, x64_c, x65_c, x68, x71_c, x72_c, x74_c, x75, x76, x79_c, x80, x81, x82_c, x84, x90, x94_c, x98);
and (w969, x3_c, x5, x7_c, x8, x9, x10, x11, x13_c, x18, x20, x21_c, x22, x23_c, x24, x27_c, x28, x29_c, x31, x33_c, x36, x37_c, x41, x42_c, x46, x49_c, x50, x51, x56_c, x58, x59, x60, x61, x64, x67, x68, x69, x71, x72, x74_c, x75, x77, x78_c, x79, x81, x86_c, x87_c, x89_c, x91, x95, x96_c, x97);
and (w970, x3_c, x6_c, x7_c, x15_c, x21, x27_c, x29_c, x32_c, x34, x36, x37, x41, x42, x48_c, x57_c, x66_c, x68, x76, x77_c, x78_c, x83_c, x93_c, x98);
and (w971, x0, x4, x5, x9, x10, x12, x17, x18_c, x19, x20, x22, x25, x26_c, x28, x29_c, x30, x32, x33_c, x34_c, x35_c, x37, x38, x39_c, x40_c, x42, x43_c, x44, x45, x47, x49, x50_c, x51, x52_c, x54, x57_c, x58_c, x59, x61_c, x62_c, x63, x65, x66, x67_c, x68_c, x69, x70, x71, x72_c, x73_c, x74_c, x76_c, x77_c, x78_c, x79_c, x80_c, x81, x82_c, x83_c, x84_c, x85_c, x87, x88_c, x89_c, x91, x92, x93_c, x95, x97, x98_c, x99);
and (w972, x0_c, x1, x2, x3, x4, x5_c, x6_c, x7_c, x8_c, x9_c, x10_c, x11_c, x12, x13, x14, x15_c, x16_c, x17_c, x18, x19, x20_c, x21, x22_c, x23_c, x24, x25_c, x26, x27, x28_c, x29_c, x32, x34_c, x35, x36, x38_c, x39, x40_c, x41_c, x42, x43_c, x44, x45, x46_c, x47, x48_c, x49_c, x50_c, x51, x52, x53, x54, x55, x56_c, x57_c, x58_c, x59, x60_c, x61, x62, x63_c, x64_c, x65_c, x66, x67, x68, x69, x70, x71_c, x72, x75_c, x76_c, x77_c, x78, x79_c, x80_c, x81_c, x82_c, x83, x84, x85_c, x86_c, x87_c, x88, x89_c, x90_c, x91_c, x92, x93, x94, x96, x98, x99);
and (w973, x0_c, x1, x2_c, x3, x4_c, x5, x6, x7_c, x8, x9, x10, x11_c, x12, x13_c, x14_c, x15, x16_c, x18_c, x19_c, x20_c, x21_c, x22, x23_c, x24_c, x25_c, x26, x27, x28, x29_c, x30_c, x31_c, x32, x33, x34_c, x35, x36_c, x37_c, x38, x39_c, x40, x41_c, x42, x43, x44_c, x45, x46, x47_c, x48, x49, x50, x51_c, x52_c, x53, x54, x55, x56_c, x57_c, x58, x59_c, x60_c, x61_c, x62, x63, x66, x67_c, x68, x69_c, x70, x71, x72, x74, x75_c, x76, x78, x79_c, x80, x82_c, x84, x85_c, x86_c, x87, x88, x89, x90_c, x91, x92, x93, x94, x95, x96_c, x97_c, x98_c);
and (w974, x0_c, x1_c, x2_c, x3_c, x4_c, x5_c, x6, x7, x8, x9, x10, x11, x12_c, x13_c, x14, x15_c, x16, x17_c, x18_c, x19, x20, x21_c, x22, x23, x24_c, x25, x26, x27, x28, x29_c, x30_c, x31, x32_c, x33, x34_c, x35, x36_c, x37, x38, x39, x40, x41_c, x42_c, x43_c, x44_c, x45_c, x46_c, x47_c, x48, x49, x50, x51, x52_c, x53_c, x54, x55_c, x56, x57, x58_c, x59_c, x60, x61, x62_c, x63, x64, x65, x66, x67, x68_c, x69_c, x70_c, x71, x72_c, x73, x74, x75, x76_c, x77, x78, x79_c, x80_c, x81_c, x82_c, x83_c, x84_c, x85, x86_c, x87, x88_c, x89, x90, x91, x92, x93_c, x94, x95, x96_c, x97_c, x98_c, x99_c);
and (w975, x9, x10_c, x16_c, x20_c, x44, x47, x52, x60_c, x76, x84_c);
and (w976, x1_c, x2, x6, x11, x12_c, x13_c, x20, x21, x30_c, x32, x37, x42, x49_c, x50_c, x52, x54, x55_c, x65_c, x71, x78, x81, x82_c, x84, x88_c, x94_c, x96_c, x97, x98_c);
and (w977, x5, x12_c, x16, x31, x44, x52, x53, x61, x73_c, x74, x75_c, x77, x78_c, x81, x82_c, x84, x87, x90);
and (w978, x18, x20_c, x34_c, x51, x58, x75_c, x82, x83_c);
and (w979, x1, x2_c, x4_c, x5_c, x7_c, x8, x9, x11_c, x12, x13_c, x16_c, x18, x20_c, x21_c, x22, x23, x24, x27_c, x29, x31, x32_c, x33, x36_c, x37, x38_c, x39, x40, x41, x42, x44, x45, x46, x47_c, x48_c, x49_c, x53_c, x54_c, x55_c, x57_c, x58, x61_c, x63, x64_c, x65, x66_c, x67_c, x68, x69_c, x70_c, x71, x72, x73, x75_c, x76_c, x77_c, x78_c, x79, x81_c, x83_c, x84_c, x88_c, x90, x91_c, x92_c, x94_c, x95_c, x98_c, x99);
and (w980, x0_c, x2, x3, x4, x5_c, x6, x7_c, x8, x9_c, x10, x11_c, x13, x14, x15_c, x16, x17_c, x18, x19_c, x20_c, x21, x22, x23, x24_c, x25, x26_c, x28, x29_c, x30_c, x31_c, x32_c, x33_c, x34, x36, x37_c, x38, x39_c, x40_c, x41, x42_c, x43, x44, x45_c, x46, x47_c, x48_c, x49_c, x50, x51, x52, x53, x54_c, x55, x56, x59, x60, x63, x64, x65, x66, x67_c, x68_c, x69, x70_c, x71_c, x72_c, x73_c, x74_c, x75, x76, x77_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x84_c, x85_c, x86, x87_c, x88, x89_c, x90_c, x94_c, x95, x96, x97_c, x98, x99);
and (w981, x1, x4, x5_c, x13_c, x15, x23, x24_c, x31, x33, x39_c, x43, x46, x49_c, x50_c, x54_c, x60_c, x67, x71_c, x74_c, x78_c, x83_c, x86_c, x87, x89_c, x93, x95_c);
and (w982, x0_c, x1_c, x2_c, x3_c, x4_c, x6, x7_c, x8_c, x9, x10, x11_c, x12, x13_c, x14_c, x15_c, x16_c, x17, x18, x19, x20, x21_c, x22, x23, x24, x25_c, x26, x27_c, x28, x29_c, x30, x31, x32_c, x33_c, x34, x35, x36_c, x37, x38_c, x39_c, x40, x41, x42_c, x43_c, x44, x45_c, x46, x47, x48_c, x49, x50_c, x51_c, x52, x53_c, x54_c, x55_c, x56, x57_c, x58, x59, x60_c, x61, x62_c, x63, x64, x65, x66_c, x67_c, x68, x69, x70_c, x71_c, x72_c, x73, x74_c, x75_c, x76, x77, x78, x79, x80_c, x81_c, x82, x83_c, x84, x85, x86, x87_c, x88_c, x89_c, x90_c, x91, x92_c, x93_c, x94, x95_c, x96, x97_c, x98_c, x99_c);
and (w983, x0_c, x1, x4_c, x5_c, x6_c, x9_c, x13, x18, x19_c, x24_c, x26, x27_c, x28_c, x29_c, x34_c, x35_c, x36_c, x38, x39, x42, x43_c, x44, x45, x46, x47, x49_c, x54, x56_c, x58, x59_c, x60, x61_c, x63, x64_c, x65_c, x66_c, x71, x73_c, x74_c, x75, x77_c, x78_c, x79, x81_c, x82, x84_c, x86_c, x87, x88_c, x89_c, x91, x93_c, x94_c, x95_c, x96_c, x98);
and (w984, x2_c, x6_c, x9, x10, x11_c, x14, x15, x16, x18, x19, x22, x24_c, x25, x26_c, x27, x28_c, x29, x30, x33_c, x34_c, x35, x36_c, x39_c, x41_c, x42_c, x43, x44, x46, x47_c, x49_c, x50, x52, x54, x55_c, x57, x60, x62, x63, x64, x65_c, x66, x67, x68, x70, x71, x72, x74_c, x75_c, x76, x77, x79, x80, x81, x83, x86, x88, x89_c, x92, x93_c, x94, x95_c, x96_c, x98);
and (w985, x0_c, x1_c, x3, x4_c, x5_c, x6, x7, x8, x10_c, x11_c, x12, x13_c, x14, x16_c, x17, x18_c, x20_c, x21_c, x22_c, x23_c, x24, x25, x26_c, x27, x28, x29, x31, x32, x33, x35_c, x37, x38, x40_c, x42_c, x43_c, x44_c, x45_c, x46, x48, x52, x56_c, x58, x59, x60, x61, x62, x63, x64, x65, x66_c, x67_c, x69_c, x70, x71, x72, x73, x74, x75, x76_c, x78_c, x79_c, x81_c, x82, x83, x84, x85_c, x86, x88_c, x89_c, x90_c, x92_c, x93, x96_c, x97_c, x99);
and (w986, x0_c, x2, x7, x9, x14, x22, x26, x28_c, x40, x54, x58, x59_c, x60, x62_c, x65_c, x70, x84_c, x98);
and (w987, x0_c, x1_c, x2_c, x4_c, x5_c, x6_c, x7_c, x8, x9, x10, x11, x12, x13, x14, x15, x18, x23, x24, x25_c, x26_c, x27_c, x28, x29_c, x31, x32_c, x33_c, x34, x35, x39, x40_c, x42_c, x44, x45_c, x47, x49_c, x50, x53_c, x54, x55_c, x57, x58, x59_c, x60, x62_c, x63_c, x67_c, x68, x70, x71_c, x73, x74_c, x76, x77, x78, x80_c, x81, x86, x87_c, x88_c, x89_c, x90, x91, x93_c, x95, x96, x97_c, x98);
and (w988, x1_c, x3, x5, x6, x9, x13, x19_c, x20_c, x28_c, x31_c, x32_c, x35, x40, x41, x43_c, x46, x48, x51_c, x55_c, x56, x57_c, x61_c, x63, x64, x65_c, x66, x67, x68, x70, x71_c, x72_c, x73_c, x74, x77_c, x87_c, x89, x90, x91_c, x97_c, x98, x99_c);
and (w989, x4_c, x10, x15_c, x22_c, x24_c, x27, x30, x34_c, x36_c, x38, x39_c, x47, x53, x54_c, x69, x71_c, x72_c, x73, x75, x81_c, x87, x90, x95_c, x97);
and (w990, x0, x1_c, x2_c, x3_c, x4_c, x5_c, x6_c, x7, x11_c, x12, x14_c, x15, x17_c, x18_c, x19_c, x20, x21, x22, x23_c, x24, x25, x26, x27, x28_c, x29, x30_c, x31, x32, x33_c, x34_c, x35_c, x36, x37, x38, x40, x41_c, x42, x43_c, x44, x45, x46, x47, x48, x49_c, x50_c, x51, x52, x53_c, x54, x55_c, x56_c, x57_c, x60, x61, x62_c, x63, x65, x66_c, x68, x69_c, x70_c, x71, x72, x73_c, x74, x76_c, x78_c, x79_c, x80, x81_c, x82_c, x83_c, x85, x86_c, x88, x89, x90, x91, x92, x93, x94, x95, x96_c, x97_c, x98_c);
and (w991, x1, x2, x3, x4, x5, x6, x7, x8_c, x9_c, x10, x12, x13, x14_c, x15, x17_c, x18, x19, x20, x21_c, x22_c, x23, x24, x25_c, x26_c, x28_c, x29_c, x30, x31, x32, x33, x36, x39, x40_c, x41_c, x42_c, x43_c, x44, x45, x46, x47, x49_c, x51, x52_c, x53, x54, x55_c, x56_c, x57_c, x58_c, x59, x60, x61_c, x62, x63_c, x64, x65_c, x66_c, x67, x68, x69, x70, x71, x72_c, x73, x76_c, x77_c, x78_c, x79, x80_c, x82_c, x84, x85_c, x87, x88_c, x89_c, x90_c, x91_c, x92_c, x93, x94, x95, x96, x97, x98_c, x99);
and (w992, x0_c, x2, x3, x4_c, x7, x8, x11, x15_c, x16_c, x17_c, x18, x22, x24, x26_c, x28_c, x30, x31_c, x32, x34_c, x35_c, x36, x37, x38_c, x40, x41, x42_c, x44, x45, x46, x47, x48, x49_c, x53_c, x54, x56_c, x57, x58_c, x60, x61, x62_c, x63, x64, x65_c, x66_c, x67_c, x68_c, x70_c, x72_c, x73, x75, x76_c, x77, x78, x81_c, x82, x83, x85_c, x88, x90, x91, x94_c, x95_c, x96_c, x97_c, x98_c, x99);
and (w993, x1_c, x4_c, x13_c, x14_c, x15, x33, x35, x38_c, x39_c, x40, x41, x46, x48, x50, x51_c, x52, x54, x56, x57_c, x58, x63_c, x64, x68, x70, x71, x72, x76, x78_c, x86_c, x88_c, x96, x99);
and (w994, x0_c, x1, x2, x3_c, x4_c, x5, x6_c, x7_c, x8, x9_c, x10_c, x11_c, x13, x14_c, x15_c, x17, x18, x19_c, x20_c, x21, x22, x23_c, x24_c, x25, x26, x27, x28, x29_c, x30_c, x31, x32_c, x33, x34, x35, x36, x37_c, x38_c, x39_c, x40, x41, x42, x43, x45_c, x46, x47, x48, x49, x50, x51, x52, x53, x54_c, x55_c, x56, x57, x59_c, x60_c, x61, x62, x63, x64_c, x65, x66, x67_c, x69_c, x70_c, x71, x72_c, x74_c, x75_c, x76_c, x77_c, x78_c, x79, x80, x81_c, x82, x84_c, x85_c, x86, x87_c, x88_c, x89, x90, x91_c, x92_c, x93_c, x94, x95, x96_c, x97, x98_c, x99_c);
and (w995, x4_c, x9_c, x11_c, x12, x25, x27, x50, x56, x58_c, x71, x81_c, x88_c, x93_c, x95_c);
and (w996, x1_c, x2_c, x6, x8, x9_c, x10_c, x12_c, x14, x16_c, x17, x18_c, x19, x20, x21_c, x22_c, x24_c, x25, x26, x30, x31_c, x34, x35_c, x36_c, x37_c, x39, x41_c, x45_c, x46_c, x50, x51, x52_c, x61, x63, x64_c, x66, x68, x69_c, x71, x72, x75, x76_c, x78, x79, x80_c, x82, x84_c, x85, x88_c, x89_c, x94_c, x96, x97, x98_c, x99_c);
and (w997, x1_c, x8_c, x19_c, x20, x29_c, x36_c, x51, x52, x54_c, x55_c, x63, x66_c, x68, x74_c, x84, x86_c, x88_c, x94_c);
and (w998, x0, x1, x2_c, x3, x4, x5_c, x6_c, x8_c, x10_c, x12, x13_c, x14, x15, x16_c, x17, x19_c, x20, x21_c, x22_c, x23_c, x24, x25_c, x26, x27_c, x28_c, x29_c, x30_c, x31_c, x32_c, x33, x34, x35_c, x37_c, x38, x40, x41, x42_c, x43, x44_c, x46_c, x48, x49_c, x50, x51_c, x52, x53_c, x55, x56, x57, x59, x60_c, x61_c, x62_c, x63, x64_c, x65_c, x66_c, x68_c, x69_c, x70_c, x71_c, x72, x73_c, x74_c, x75, x76_c, x78, x79, x80, x81_c, x82_c, x83_c, x84_c, x86, x87, x88_c, x90_c, x92_c, x95, x96, x97_c, x99_c);
and (w999, x4, x6_c, x7, x8, x9, x10, x18, x25, x28, x31_c, x34, x36, x37_c, x38, x40, x41_c, x42_c, x43_c, x45, x46_c, x56_c, x58_c, x60, x62, x64, x69_c, x71, x72_c, x73_c, x77, x78, x81_c, x83, x85, x89_c, x90_c, x93, x94_c, x96, x99);
xor (o, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999);
endmodule
